module cc_dir_ext(
  input  [9:0]   RW0_addr,
  input          RW0_clk,
  input  [127:0] RW0_wdata,
  output [127:0] RW0_rdata,
  input          RW0_en,
  input          RW0_wmode,
  input  [7:0]   RW0_wmask
);
  wire [9:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [15:0] mem_0_0_RW0_wdata;
  wire [15:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [9:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [15:0] mem_0_1_RW0_wdata;
  wire [15:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [9:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [15:0] mem_0_2_RW0_wdata;
  wire [15:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [9:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [15:0] mem_0_3_RW0_wdata;
  wire [15:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [9:0] mem_0_4_RW0_addr;
  wire  mem_0_4_RW0_clk;
  wire [15:0] mem_0_4_RW0_wdata;
  wire [15:0] mem_0_4_RW0_rdata;
  wire  mem_0_4_RW0_en;
  wire  mem_0_4_RW0_wmode;
  wire  mem_0_4_RW0_wmask;
  wire [9:0] mem_0_5_RW0_addr;
  wire  mem_0_5_RW0_clk;
  wire [15:0] mem_0_5_RW0_wdata;
  wire [15:0] mem_0_5_RW0_rdata;
  wire  mem_0_5_RW0_en;
  wire  mem_0_5_RW0_wmode;
  wire  mem_0_5_RW0_wmask;
  wire [9:0] mem_0_6_RW0_addr;
  wire  mem_0_6_RW0_clk;
  wire [15:0] mem_0_6_RW0_wdata;
  wire [15:0] mem_0_6_RW0_rdata;
  wire  mem_0_6_RW0_en;
  wire  mem_0_6_RW0_wmode;
  wire  mem_0_6_RW0_wmask;
  wire [9:0] mem_0_7_RW0_addr;
  wire  mem_0_7_RW0_clk;
  wire [15:0] mem_0_7_RW0_wdata;
  wire [15:0] mem_0_7_RW0_rdata;
  wire  mem_0_7_RW0_en;
  wire  mem_0_7_RW0_wmode;
  wire  mem_0_7_RW0_wmask;
  wire [15:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [15:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [15:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [15:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [15:0] RW0_rdata_0_4 = mem_0_4_RW0_rdata;
  wire [15:0] RW0_rdata_0_5 = mem_0_5_RW0_rdata;
  wire [15:0] RW0_rdata_0_6 = mem_0_6_RW0_rdata;
  wire [15:0] RW0_rdata_0_7 = mem_0_7_RW0_rdata;
  wire [31:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [47:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [63:0] _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [79:0] _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [95:0] _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [111:0] _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  wire [127:0] RW0_rdata_0 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0};
  wire [31:0] _GEN_6 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [47:0] _GEN_7 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [63:0] _GEN_8 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [79:0] _GEN_9 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [95:0] _GEN_10 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [111:0] _GEN_11 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  split_cc_dir_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_cc_dir_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_cc_dir_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_cc_dir_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_cc_dir_ext mem_0_4 (
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_cc_dir_ext mem_0_5 (
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_cc_dir_ext mem_0_6 (
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_cc_dir_ext mem_0_7 (
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_7,_GEN_5};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[15:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[31:16];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[47:32];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[63:48];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
  assign mem_0_4_RW0_addr = RW0_addr;
  assign mem_0_4_RW0_clk = RW0_clk;
  assign mem_0_4_RW0_wdata = RW0_wdata[79:64];
  assign mem_0_4_RW0_en = RW0_en;
  assign mem_0_4_RW0_wmode = RW0_wmode;
  assign mem_0_4_RW0_wmask = RW0_wmask[4];
  assign mem_0_5_RW0_addr = RW0_addr;
  assign mem_0_5_RW0_clk = RW0_clk;
  assign mem_0_5_RW0_wdata = RW0_wdata[95:80];
  assign mem_0_5_RW0_en = RW0_en;
  assign mem_0_5_RW0_wmode = RW0_wmode;
  assign mem_0_5_RW0_wmask = RW0_wmask[5];
  assign mem_0_6_RW0_addr = RW0_addr;
  assign mem_0_6_RW0_clk = RW0_clk;
  assign mem_0_6_RW0_wdata = RW0_wdata[111:96];
  assign mem_0_6_RW0_en = RW0_en;
  assign mem_0_6_RW0_wmode = RW0_wmode;
  assign mem_0_6_RW0_wmask = RW0_wmask[6];
  assign mem_0_7_RW0_addr = RW0_addr;
  assign mem_0_7_RW0_clk = RW0_clk;
  assign mem_0_7_RW0_wdata = RW0_wdata[127:112];
  assign mem_0_7_RW0_en = RW0_en;
  assign mem_0_7_RW0_wmode = RW0_wmode;
  assign mem_0_7_RW0_wmask = RW0_wmask[7];
endmodule
module cc_banks_0_ext(
  input  [12:0] RW0_addr,
  input         RW0_clk,
  input  [63:0] RW0_wdata,
  output [63:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
  wire [12:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [63:0] mem_0_0_RW0_wdata;
  wire [63:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire [63:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [63:0] RW0_rdata_0 = RW0_rdata_0_0;
  split_cc_banks_0_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata = mem_0_0_RW0_rdata;
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata;
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
endmodule
module data_arrays_0_ext(
  input  [7:0]   RW0_addr,
  input          RW0_clk,
  input  [255:0] RW0_wdata,
  output [255:0] RW0_rdata,
  input          RW0_en,
  input          RW0_wmode,
  input  [31:0]  RW0_wmask
);
  wire [7:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [7:0] mem_0_0_RW0_wdata;
  wire [7:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [7:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [7:0] mem_0_1_RW0_wdata;
  wire [7:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [7:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [7:0] mem_0_2_RW0_wdata;
  wire [7:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [7:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [7:0] mem_0_3_RW0_wdata;
  wire [7:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [7:0] mem_0_4_RW0_addr;
  wire  mem_0_4_RW0_clk;
  wire [7:0] mem_0_4_RW0_wdata;
  wire [7:0] mem_0_4_RW0_rdata;
  wire  mem_0_4_RW0_en;
  wire  mem_0_4_RW0_wmode;
  wire  mem_0_4_RW0_wmask;
  wire [7:0] mem_0_5_RW0_addr;
  wire  mem_0_5_RW0_clk;
  wire [7:0] mem_0_5_RW0_wdata;
  wire [7:0] mem_0_5_RW0_rdata;
  wire  mem_0_5_RW0_en;
  wire  mem_0_5_RW0_wmode;
  wire  mem_0_5_RW0_wmask;
  wire [7:0] mem_0_6_RW0_addr;
  wire  mem_0_6_RW0_clk;
  wire [7:0] mem_0_6_RW0_wdata;
  wire [7:0] mem_0_6_RW0_rdata;
  wire  mem_0_6_RW0_en;
  wire  mem_0_6_RW0_wmode;
  wire  mem_0_6_RW0_wmask;
  wire [7:0] mem_0_7_RW0_addr;
  wire  mem_0_7_RW0_clk;
  wire [7:0] mem_0_7_RW0_wdata;
  wire [7:0] mem_0_7_RW0_rdata;
  wire  mem_0_7_RW0_en;
  wire  mem_0_7_RW0_wmode;
  wire  mem_0_7_RW0_wmask;
  wire [7:0] mem_0_8_RW0_addr;
  wire  mem_0_8_RW0_clk;
  wire [7:0] mem_0_8_RW0_wdata;
  wire [7:0] mem_0_8_RW0_rdata;
  wire  mem_0_8_RW0_en;
  wire  mem_0_8_RW0_wmode;
  wire  mem_0_8_RW0_wmask;
  wire [7:0] mem_0_9_RW0_addr;
  wire  mem_0_9_RW0_clk;
  wire [7:0] mem_0_9_RW0_wdata;
  wire [7:0] mem_0_9_RW0_rdata;
  wire  mem_0_9_RW0_en;
  wire  mem_0_9_RW0_wmode;
  wire  mem_0_9_RW0_wmask;
  wire [7:0] mem_0_10_RW0_addr;
  wire  mem_0_10_RW0_clk;
  wire [7:0] mem_0_10_RW0_wdata;
  wire [7:0] mem_0_10_RW0_rdata;
  wire  mem_0_10_RW0_en;
  wire  mem_0_10_RW0_wmode;
  wire  mem_0_10_RW0_wmask;
  wire [7:0] mem_0_11_RW0_addr;
  wire  mem_0_11_RW0_clk;
  wire [7:0] mem_0_11_RW0_wdata;
  wire [7:0] mem_0_11_RW0_rdata;
  wire  mem_0_11_RW0_en;
  wire  mem_0_11_RW0_wmode;
  wire  mem_0_11_RW0_wmask;
  wire [7:0] mem_0_12_RW0_addr;
  wire  mem_0_12_RW0_clk;
  wire [7:0] mem_0_12_RW0_wdata;
  wire [7:0] mem_0_12_RW0_rdata;
  wire  mem_0_12_RW0_en;
  wire  mem_0_12_RW0_wmode;
  wire  mem_0_12_RW0_wmask;
  wire [7:0] mem_0_13_RW0_addr;
  wire  mem_0_13_RW0_clk;
  wire [7:0] mem_0_13_RW0_wdata;
  wire [7:0] mem_0_13_RW0_rdata;
  wire  mem_0_13_RW0_en;
  wire  mem_0_13_RW0_wmode;
  wire  mem_0_13_RW0_wmask;
  wire [7:0] mem_0_14_RW0_addr;
  wire  mem_0_14_RW0_clk;
  wire [7:0] mem_0_14_RW0_wdata;
  wire [7:0] mem_0_14_RW0_rdata;
  wire  mem_0_14_RW0_en;
  wire  mem_0_14_RW0_wmode;
  wire  mem_0_14_RW0_wmask;
  wire [7:0] mem_0_15_RW0_addr;
  wire  mem_0_15_RW0_clk;
  wire [7:0] mem_0_15_RW0_wdata;
  wire [7:0] mem_0_15_RW0_rdata;
  wire  mem_0_15_RW0_en;
  wire  mem_0_15_RW0_wmode;
  wire  mem_0_15_RW0_wmask;
  wire [7:0] mem_0_16_RW0_addr;
  wire  mem_0_16_RW0_clk;
  wire [7:0] mem_0_16_RW0_wdata;
  wire [7:0] mem_0_16_RW0_rdata;
  wire  mem_0_16_RW0_en;
  wire  mem_0_16_RW0_wmode;
  wire  mem_0_16_RW0_wmask;
  wire [7:0] mem_0_17_RW0_addr;
  wire  mem_0_17_RW0_clk;
  wire [7:0] mem_0_17_RW0_wdata;
  wire [7:0] mem_0_17_RW0_rdata;
  wire  mem_0_17_RW0_en;
  wire  mem_0_17_RW0_wmode;
  wire  mem_0_17_RW0_wmask;
  wire [7:0] mem_0_18_RW0_addr;
  wire  mem_0_18_RW0_clk;
  wire [7:0] mem_0_18_RW0_wdata;
  wire [7:0] mem_0_18_RW0_rdata;
  wire  mem_0_18_RW0_en;
  wire  mem_0_18_RW0_wmode;
  wire  mem_0_18_RW0_wmask;
  wire [7:0] mem_0_19_RW0_addr;
  wire  mem_0_19_RW0_clk;
  wire [7:0] mem_0_19_RW0_wdata;
  wire [7:0] mem_0_19_RW0_rdata;
  wire  mem_0_19_RW0_en;
  wire  mem_0_19_RW0_wmode;
  wire  mem_0_19_RW0_wmask;
  wire [7:0] mem_0_20_RW0_addr;
  wire  mem_0_20_RW0_clk;
  wire [7:0] mem_0_20_RW0_wdata;
  wire [7:0] mem_0_20_RW0_rdata;
  wire  mem_0_20_RW0_en;
  wire  mem_0_20_RW0_wmode;
  wire  mem_0_20_RW0_wmask;
  wire [7:0] mem_0_21_RW0_addr;
  wire  mem_0_21_RW0_clk;
  wire [7:0] mem_0_21_RW0_wdata;
  wire [7:0] mem_0_21_RW0_rdata;
  wire  mem_0_21_RW0_en;
  wire  mem_0_21_RW0_wmode;
  wire  mem_0_21_RW0_wmask;
  wire [7:0] mem_0_22_RW0_addr;
  wire  mem_0_22_RW0_clk;
  wire [7:0] mem_0_22_RW0_wdata;
  wire [7:0] mem_0_22_RW0_rdata;
  wire  mem_0_22_RW0_en;
  wire  mem_0_22_RW0_wmode;
  wire  mem_0_22_RW0_wmask;
  wire [7:0] mem_0_23_RW0_addr;
  wire  mem_0_23_RW0_clk;
  wire [7:0] mem_0_23_RW0_wdata;
  wire [7:0] mem_0_23_RW0_rdata;
  wire  mem_0_23_RW0_en;
  wire  mem_0_23_RW0_wmode;
  wire  mem_0_23_RW0_wmask;
  wire [7:0] mem_0_24_RW0_addr;
  wire  mem_0_24_RW0_clk;
  wire [7:0] mem_0_24_RW0_wdata;
  wire [7:0] mem_0_24_RW0_rdata;
  wire  mem_0_24_RW0_en;
  wire  mem_0_24_RW0_wmode;
  wire  mem_0_24_RW0_wmask;
  wire [7:0] mem_0_25_RW0_addr;
  wire  mem_0_25_RW0_clk;
  wire [7:0] mem_0_25_RW0_wdata;
  wire [7:0] mem_0_25_RW0_rdata;
  wire  mem_0_25_RW0_en;
  wire  mem_0_25_RW0_wmode;
  wire  mem_0_25_RW0_wmask;
  wire [7:0] mem_0_26_RW0_addr;
  wire  mem_0_26_RW0_clk;
  wire [7:0] mem_0_26_RW0_wdata;
  wire [7:0] mem_0_26_RW0_rdata;
  wire  mem_0_26_RW0_en;
  wire  mem_0_26_RW0_wmode;
  wire  mem_0_26_RW0_wmask;
  wire [7:0] mem_0_27_RW0_addr;
  wire  mem_0_27_RW0_clk;
  wire [7:0] mem_0_27_RW0_wdata;
  wire [7:0] mem_0_27_RW0_rdata;
  wire  mem_0_27_RW0_en;
  wire  mem_0_27_RW0_wmode;
  wire  mem_0_27_RW0_wmask;
  wire [7:0] mem_0_28_RW0_addr;
  wire  mem_0_28_RW0_clk;
  wire [7:0] mem_0_28_RW0_wdata;
  wire [7:0] mem_0_28_RW0_rdata;
  wire  mem_0_28_RW0_en;
  wire  mem_0_28_RW0_wmode;
  wire  mem_0_28_RW0_wmask;
  wire [7:0] mem_0_29_RW0_addr;
  wire  mem_0_29_RW0_clk;
  wire [7:0] mem_0_29_RW0_wdata;
  wire [7:0] mem_0_29_RW0_rdata;
  wire  mem_0_29_RW0_en;
  wire  mem_0_29_RW0_wmode;
  wire  mem_0_29_RW0_wmask;
  wire [7:0] mem_0_30_RW0_addr;
  wire  mem_0_30_RW0_clk;
  wire [7:0] mem_0_30_RW0_wdata;
  wire [7:0] mem_0_30_RW0_rdata;
  wire  mem_0_30_RW0_en;
  wire  mem_0_30_RW0_wmode;
  wire  mem_0_30_RW0_wmask;
  wire [7:0] mem_0_31_RW0_addr;
  wire  mem_0_31_RW0_clk;
  wire [7:0] mem_0_31_RW0_wdata;
  wire [7:0] mem_0_31_RW0_rdata;
  wire  mem_0_31_RW0_en;
  wire  mem_0_31_RW0_wmode;
  wire  mem_0_31_RW0_wmask;
  wire [7:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [7:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [7:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [7:0] RW0_rdata_0_4 = mem_0_4_RW0_rdata;
  wire [7:0] RW0_rdata_0_5 = mem_0_5_RW0_rdata;
  wire [7:0] RW0_rdata_0_6 = mem_0_6_RW0_rdata;
  wire [7:0] RW0_rdata_0_7 = mem_0_7_RW0_rdata;
  wire [7:0] RW0_rdata_0_8 = mem_0_8_RW0_rdata;
  wire [7:0] RW0_rdata_0_9 = mem_0_9_RW0_rdata;
  wire [7:0] RW0_rdata_0_10 = mem_0_10_RW0_rdata;
  wire [7:0] RW0_rdata_0_11 = mem_0_11_RW0_rdata;
  wire [7:0] RW0_rdata_0_12 = mem_0_12_RW0_rdata;
  wire [7:0] RW0_rdata_0_13 = mem_0_13_RW0_rdata;
  wire [7:0] RW0_rdata_0_14 = mem_0_14_RW0_rdata;
  wire [7:0] RW0_rdata_0_15 = mem_0_15_RW0_rdata;
  wire [7:0] RW0_rdata_0_16 = mem_0_16_RW0_rdata;
  wire [7:0] RW0_rdata_0_17 = mem_0_17_RW0_rdata;
  wire [7:0] RW0_rdata_0_18 = mem_0_18_RW0_rdata;
  wire [7:0] RW0_rdata_0_19 = mem_0_19_RW0_rdata;
  wire [7:0] RW0_rdata_0_20 = mem_0_20_RW0_rdata;
  wire [7:0] RW0_rdata_0_21 = mem_0_21_RW0_rdata;
  wire [7:0] RW0_rdata_0_22 = mem_0_22_RW0_rdata;
  wire [7:0] RW0_rdata_0_23 = mem_0_23_RW0_rdata;
  wire [7:0] RW0_rdata_0_24 = mem_0_24_RW0_rdata;
  wire [7:0] RW0_rdata_0_25 = mem_0_25_RW0_rdata;
  wire [7:0] RW0_rdata_0_26 = mem_0_26_RW0_rdata;
  wire [7:0] RW0_rdata_0_27 = mem_0_27_RW0_rdata;
  wire [7:0] RW0_rdata_0_28 = mem_0_28_RW0_rdata;
  wire [7:0] RW0_rdata_0_29 = mem_0_29_RW0_rdata;
  wire [7:0] RW0_rdata_0_30 = mem_0_30_RW0_rdata;
  wire [7:0] RW0_rdata_0_31 = mem_0_31_RW0_rdata;
  wire [15:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [31:0] _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [39:0] _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [47:0] _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [55:0] _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  wire [63:0] _GEN_6 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0};
  wire [71:0] _GEN_7 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,
    RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [79:0] _GEN_8 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,
    RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [87:0] _GEN_9 = {RW0_rdata_0_10,_GEN_8};
  wire [95:0] _GEN_10 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [103:0] _GEN_11 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [111:0] _GEN_12 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [119:0] _GEN_13 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [127:0] _GEN_14 = {RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,
    _GEN_8};
  wire [135:0] _GEN_15 = {RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,
    RW0_rdata_0_10,_GEN_8};
  wire [143:0] _GEN_16 = {RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,
    RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [151:0] _GEN_17 = {RW0_rdata_0_18,RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,
    RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [159:0] _GEN_18 = {RW0_rdata_0_19,_GEN_17};
  wire [167:0] _GEN_19 = {RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [175:0] _GEN_20 = {RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [183:0] _GEN_21 = {RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [191:0] _GEN_22 = {RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [199:0] _GEN_23 = {RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,
    _GEN_17};
  wire [207:0] _GEN_24 = {RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,
    RW0_rdata_0_19,_GEN_17};
  wire [215:0] _GEN_25 = {RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,
    RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [223:0] _GEN_26 = {RW0_rdata_0_27,RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,
    RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [231:0] _GEN_27 = {RW0_rdata_0_28,_GEN_26};
  wire [239:0] _GEN_28 = {RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  wire [247:0] _GEN_29 = {RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  wire [255:0] RW0_rdata_0 = {RW0_rdata_0_31,RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  wire [15:0] _GEN_30 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_31 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [31:0] _GEN_32 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [39:0] _GEN_33 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [47:0] _GEN_34 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [55:0] _GEN_35 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  wire [63:0] _GEN_36 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0};
  wire [71:0] _GEN_37 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,
    RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [79:0] _GEN_38 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,
    RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [87:0] _GEN_39 = {RW0_rdata_0_10,_GEN_8};
  wire [95:0] _GEN_40 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [103:0] _GEN_41 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [111:0] _GEN_42 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [119:0] _GEN_43 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [127:0] _GEN_44 = {RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,
    _GEN_8};
  wire [135:0] _GEN_45 = {RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,
    RW0_rdata_0_10,_GEN_8};
  wire [143:0] _GEN_46 = {RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,
    RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [151:0] _GEN_47 = {RW0_rdata_0_18,RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,
    RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [159:0] _GEN_48 = {RW0_rdata_0_19,_GEN_17};
  wire [167:0] _GEN_49 = {RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [175:0] _GEN_50 = {RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [183:0] _GEN_51 = {RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [191:0] _GEN_52 = {RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [199:0] _GEN_53 = {RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,
    _GEN_17};
  wire [207:0] _GEN_54 = {RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,
    RW0_rdata_0_19,_GEN_17};
  wire [215:0] _GEN_55 = {RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,
    RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [223:0] _GEN_56 = {RW0_rdata_0_27,RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,
    RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17};
  wire [231:0] _GEN_57 = {RW0_rdata_0_28,_GEN_26};
  wire [239:0] _GEN_58 = {RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  wire [247:0] _GEN_59 = {RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26};
  split_data_arrays_0_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_4 (
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_5 (
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_6 (
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_7 (
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_8 (
    .RW0_addr(mem_0_8_RW0_addr),
    .RW0_clk(mem_0_8_RW0_clk),
    .RW0_wdata(mem_0_8_RW0_wdata),
    .RW0_rdata(mem_0_8_RW0_rdata),
    .RW0_en(mem_0_8_RW0_en),
    .RW0_wmode(mem_0_8_RW0_wmode),
    .RW0_wmask(mem_0_8_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_9 (
    .RW0_addr(mem_0_9_RW0_addr),
    .RW0_clk(mem_0_9_RW0_clk),
    .RW0_wdata(mem_0_9_RW0_wdata),
    .RW0_rdata(mem_0_9_RW0_rdata),
    .RW0_en(mem_0_9_RW0_en),
    .RW0_wmode(mem_0_9_RW0_wmode),
    .RW0_wmask(mem_0_9_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_10 (
    .RW0_addr(mem_0_10_RW0_addr),
    .RW0_clk(mem_0_10_RW0_clk),
    .RW0_wdata(mem_0_10_RW0_wdata),
    .RW0_rdata(mem_0_10_RW0_rdata),
    .RW0_en(mem_0_10_RW0_en),
    .RW0_wmode(mem_0_10_RW0_wmode),
    .RW0_wmask(mem_0_10_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_11 (
    .RW0_addr(mem_0_11_RW0_addr),
    .RW0_clk(mem_0_11_RW0_clk),
    .RW0_wdata(mem_0_11_RW0_wdata),
    .RW0_rdata(mem_0_11_RW0_rdata),
    .RW0_en(mem_0_11_RW0_en),
    .RW0_wmode(mem_0_11_RW0_wmode),
    .RW0_wmask(mem_0_11_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_12 (
    .RW0_addr(mem_0_12_RW0_addr),
    .RW0_clk(mem_0_12_RW0_clk),
    .RW0_wdata(mem_0_12_RW0_wdata),
    .RW0_rdata(mem_0_12_RW0_rdata),
    .RW0_en(mem_0_12_RW0_en),
    .RW0_wmode(mem_0_12_RW0_wmode),
    .RW0_wmask(mem_0_12_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_13 (
    .RW0_addr(mem_0_13_RW0_addr),
    .RW0_clk(mem_0_13_RW0_clk),
    .RW0_wdata(mem_0_13_RW0_wdata),
    .RW0_rdata(mem_0_13_RW0_rdata),
    .RW0_en(mem_0_13_RW0_en),
    .RW0_wmode(mem_0_13_RW0_wmode),
    .RW0_wmask(mem_0_13_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_14 (
    .RW0_addr(mem_0_14_RW0_addr),
    .RW0_clk(mem_0_14_RW0_clk),
    .RW0_wdata(mem_0_14_RW0_wdata),
    .RW0_rdata(mem_0_14_RW0_rdata),
    .RW0_en(mem_0_14_RW0_en),
    .RW0_wmode(mem_0_14_RW0_wmode),
    .RW0_wmask(mem_0_14_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_15 (
    .RW0_addr(mem_0_15_RW0_addr),
    .RW0_clk(mem_0_15_RW0_clk),
    .RW0_wdata(mem_0_15_RW0_wdata),
    .RW0_rdata(mem_0_15_RW0_rdata),
    .RW0_en(mem_0_15_RW0_en),
    .RW0_wmode(mem_0_15_RW0_wmode),
    .RW0_wmask(mem_0_15_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_16 (
    .RW0_addr(mem_0_16_RW0_addr),
    .RW0_clk(mem_0_16_RW0_clk),
    .RW0_wdata(mem_0_16_RW0_wdata),
    .RW0_rdata(mem_0_16_RW0_rdata),
    .RW0_en(mem_0_16_RW0_en),
    .RW0_wmode(mem_0_16_RW0_wmode),
    .RW0_wmask(mem_0_16_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_17 (
    .RW0_addr(mem_0_17_RW0_addr),
    .RW0_clk(mem_0_17_RW0_clk),
    .RW0_wdata(mem_0_17_RW0_wdata),
    .RW0_rdata(mem_0_17_RW0_rdata),
    .RW0_en(mem_0_17_RW0_en),
    .RW0_wmode(mem_0_17_RW0_wmode),
    .RW0_wmask(mem_0_17_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_18 (
    .RW0_addr(mem_0_18_RW0_addr),
    .RW0_clk(mem_0_18_RW0_clk),
    .RW0_wdata(mem_0_18_RW0_wdata),
    .RW0_rdata(mem_0_18_RW0_rdata),
    .RW0_en(mem_0_18_RW0_en),
    .RW0_wmode(mem_0_18_RW0_wmode),
    .RW0_wmask(mem_0_18_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_19 (
    .RW0_addr(mem_0_19_RW0_addr),
    .RW0_clk(mem_0_19_RW0_clk),
    .RW0_wdata(mem_0_19_RW0_wdata),
    .RW0_rdata(mem_0_19_RW0_rdata),
    .RW0_en(mem_0_19_RW0_en),
    .RW0_wmode(mem_0_19_RW0_wmode),
    .RW0_wmask(mem_0_19_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_20 (
    .RW0_addr(mem_0_20_RW0_addr),
    .RW0_clk(mem_0_20_RW0_clk),
    .RW0_wdata(mem_0_20_RW0_wdata),
    .RW0_rdata(mem_0_20_RW0_rdata),
    .RW0_en(mem_0_20_RW0_en),
    .RW0_wmode(mem_0_20_RW0_wmode),
    .RW0_wmask(mem_0_20_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_21 (
    .RW0_addr(mem_0_21_RW0_addr),
    .RW0_clk(mem_0_21_RW0_clk),
    .RW0_wdata(mem_0_21_RW0_wdata),
    .RW0_rdata(mem_0_21_RW0_rdata),
    .RW0_en(mem_0_21_RW0_en),
    .RW0_wmode(mem_0_21_RW0_wmode),
    .RW0_wmask(mem_0_21_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_22 (
    .RW0_addr(mem_0_22_RW0_addr),
    .RW0_clk(mem_0_22_RW0_clk),
    .RW0_wdata(mem_0_22_RW0_wdata),
    .RW0_rdata(mem_0_22_RW0_rdata),
    .RW0_en(mem_0_22_RW0_en),
    .RW0_wmode(mem_0_22_RW0_wmode),
    .RW0_wmask(mem_0_22_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_23 (
    .RW0_addr(mem_0_23_RW0_addr),
    .RW0_clk(mem_0_23_RW0_clk),
    .RW0_wdata(mem_0_23_RW0_wdata),
    .RW0_rdata(mem_0_23_RW0_rdata),
    .RW0_en(mem_0_23_RW0_en),
    .RW0_wmode(mem_0_23_RW0_wmode),
    .RW0_wmask(mem_0_23_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_24 (
    .RW0_addr(mem_0_24_RW0_addr),
    .RW0_clk(mem_0_24_RW0_clk),
    .RW0_wdata(mem_0_24_RW0_wdata),
    .RW0_rdata(mem_0_24_RW0_rdata),
    .RW0_en(mem_0_24_RW0_en),
    .RW0_wmode(mem_0_24_RW0_wmode),
    .RW0_wmask(mem_0_24_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_25 (
    .RW0_addr(mem_0_25_RW0_addr),
    .RW0_clk(mem_0_25_RW0_clk),
    .RW0_wdata(mem_0_25_RW0_wdata),
    .RW0_rdata(mem_0_25_RW0_rdata),
    .RW0_en(mem_0_25_RW0_en),
    .RW0_wmode(mem_0_25_RW0_wmode),
    .RW0_wmask(mem_0_25_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_26 (
    .RW0_addr(mem_0_26_RW0_addr),
    .RW0_clk(mem_0_26_RW0_clk),
    .RW0_wdata(mem_0_26_RW0_wdata),
    .RW0_rdata(mem_0_26_RW0_rdata),
    .RW0_en(mem_0_26_RW0_en),
    .RW0_wmode(mem_0_26_RW0_wmode),
    .RW0_wmask(mem_0_26_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_27 (
    .RW0_addr(mem_0_27_RW0_addr),
    .RW0_clk(mem_0_27_RW0_clk),
    .RW0_wdata(mem_0_27_RW0_wdata),
    .RW0_rdata(mem_0_27_RW0_rdata),
    .RW0_en(mem_0_27_RW0_en),
    .RW0_wmode(mem_0_27_RW0_wmode),
    .RW0_wmask(mem_0_27_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_28 (
    .RW0_addr(mem_0_28_RW0_addr),
    .RW0_clk(mem_0_28_RW0_clk),
    .RW0_wdata(mem_0_28_RW0_wdata),
    .RW0_rdata(mem_0_28_RW0_rdata),
    .RW0_en(mem_0_28_RW0_en),
    .RW0_wmode(mem_0_28_RW0_wmode),
    .RW0_wmask(mem_0_28_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_29 (
    .RW0_addr(mem_0_29_RW0_addr),
    .RW0_clk(mem_0_29_RW0_clk),
    .RW0_wdata(mem_0_29_RW0_wdata),
    .RW0_rdata(mem_0_29_RW0_rdata),
    .RW0_en(mem_0_29_RW0_en),
    .RW0_wmode(mem_0_29_RW0_wmode),
    .RW0_wmask(mem_0_29_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_30 (
    .RW0_addr(mem_0_30_RW0_addr),
    .RW0_clk(mem_0_30_RW0_clk),
    .RW0_wdata(mem_0_30_RW0_wdata),
    .RW0_rdata(mem_0_30_RW0_rdata),
    .RW0_en(mem_0_30_RW0_en),
    .RW0_wmode(mem_0_30_RW0_wmode),
    .RW0_wmask(mem_0_30_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_31 (
    .RW0_addr(mem_0_31_RW0_addr),
    .RW0_clk(mem_0_31_RW0_clk),
    .RW0_wdata(mem_0_31_RW0_wdata),
    .RW0_rdata(mem_0_31_RW0_rdata),
    .RW0_en(mem_0_31_RW0_en),
    .RW0_wmode(mem_0_31_RW0_wmode),
    .RW0_wmask(mem_0_31_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_31,_GEN_29};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[7:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[15:8];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[23:16];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[31:24];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
  assign mem_0_4_RW0_addr = RW0_addr;
  assign mem_0_4_RW0_clk = RW0_clk;
  assign mem_0_4_RW0_wdata = RW0_wdata[39:32];
  assign mem_0_4_RW0_en = RW0_en;
  assign mem_0_4_RW0_wmode = RW0_wmode;
  assign mem_0_4_RW0_wmask = RW0_wmask[4];
  assign mem_0_5_RW0_addr = RW0_addr;
  assign mem_0_5_RW0_clk = RW0_clk;
  assign mem_0_5_RW0_wdata = RW0_wdata[47:40];
  assign mem_0_5_RW0_en = RW0_en;
  assign mem_0_5_RW0_wmode = RW0_wmode;
  assign mem_0_5_RW0_wmask = RW0_wmask[5];
  assign mem_0_6_RW0_addr = RW0_addr;
  assign mem_0_6_RW0_clk = RW0_clk;
  assign mem_0_6_RW0_wdata = RW0_wdata[55:48];
  assign mem_0_6_RW0_en = RW0_en;
  assign mem_0_6_RW0_wmode = RW0_wmode;
  assign mem_0_6_RW0_wmask = RW0_wmask[6];
  assign mem_0_7_RW0_addr = RW0_addr;
  assign mem_0_7_RW0_clk = RW0_clk;
  assign mem_0_7_RW0_wdata = RW0_wdata[63:56];
  assign mem_0_7_RW0_en = RW0_en;
  assign mem_0_7_RW0_wmode = RW0_wmode;
  assign mem_0_7_RW0_wmask = RW0_wmask[7];
  assign mem_0_8_RW0_addr = RW0_addr;
  assign mem_0_8_RW0_clk = RW0_clk;
  assign mem_0_8_RW0_wdata = RW0_wdata[71:64];
  assign mem_0_8_RW0_en = RW0_en;
  assign mem_0_8_RW0_wmode = RW0_wmode;
  assign mem_0_8_RW0_wmask = RW0_wmask[8];
  assign mem_0_9_RW0_addr = RW0_addr;
  assign mem_0_9_RW0_clk = RW0_clk;
  assign mem_0_9_RW0_wdata = RW0_wdata[79:72];
  assign mem_0_9_RW0_en = RW0_en;
  assign mem_0_9_RW0_wmode = RW0_wmode;
  assign mem_0_9_RW0_wmask = RW0_wmask[9];
  assign mem_0_10_RW0_addr = RW0_addr;
  assign mem_0_10_RW0_clk = RW0_clk;
  assign mem_0_10_RW0_wdata = RW0_wdata[87:80];
  assign mem_0_10_RW0_en = RW0_en;
  assign mem_0_10_RW0_wmode = RW0_wmode;
  assign mem_0_10_RW0_wmask = RW0_wmask[10];
  assign mem_0_11_RW0_addr = RW0_addr;
  assign mem_0_11_RW0_clk = RW0_clk;
  assign mem_0_11_RW0_wdata = RW0_wdata[95:88];
  assign mem_0_11_RW0_en = RW0_en;
  assign mem_0_11_RW0_wmode = RW0_wmode;
  assign mem_0_11_RW0_wmask = RW0_wmask[11];
  assign mem_0_12_RW0_addr = RW0_addr;
  assign mem_0_12_RW0_clk = RW0_clk;
  assign mem_0_12_RW0_wdata = RW0_wdata[103:96];
  assign mem_0_12_RW0_en = RW0_en;
  assign mem_0_12_RW0_wmode = RW0_wmode;
  assign mem_0_12_RW0_wmask = RW0_wmask[12];
  assign mem_0_13_RW0_addr = RW0_addr;
  assign mem_0_13_RW0_clk = RW0_clk;
  assign mem_0_13_RW0_wdata = RW0_wdata[111:104];
  assign mem_0_13_RW0_en = RW0_en;
  assign mem_0_13_RW0_wmode = RW0_wmode;
  assign mem_0_13_RW0_wmask = RW0_wmask[13];
  assign mem_0_14_RW0_addr = RW0_addr;
  assign mem_0_14_RW0_clk = RW0_clk;
  assign mem_0_14_RW0_wdata = RW0_wdata[119:112];
  assign mem_0_14_RW0_en = RW0_en;
  assign mem_0_14_RW0_wmode = RW0_wmode;
  assign mem_0_14_RW0_wmask = RW0_wmask[14];
  assign mem_0_15_RW0_addr = RW0_addr;
  assign mem_0_15_RW0_clk = RW0_clk;
  assign mem_0_15_RW0_wdata = RW0_wdata[127:120];
  assign mem_0_15_RW0_en = RW0_en;
  assign mem_0_15_RW0_wmode = RW0_wmode;
  assign mem_0_15_RW0_wmask = RW0_wmask[15];
  assign mem_0_16_RW0_addr = RW0_addr;
  assign mem_0_16_RW0_clk = RW0_clk;
  assign mem_0_16_RW0_wdata = RW0_wdata[135:128];
  assign mem_0_16_RW0_en = RW0_en;
  assign mem_0_16_RW0_wmode = RW0_wmode;
  assign mem_0_16_RW0_wmask = RW0_wmask[16];
  assign mem_0_17_RW0_addr = RW0_addr;
  assign mem_0_17_RW0_clk = RW0_clk;
  assign mem_0_17_RW0_wdata = RW0_wdata[143:136];
  assign mem_0_17_RW0_en = RW0_en;
  assign mem_0_17_RW0_wmode = RW0_wmode;
  assign mem_0_17_RW0_wmask = RW0_wmask[17];
  assign mem_0_18_RW0_addr = RW0_addr;
  assign mem_0_18_RW0_clk = RW0_clk;
  assign mem_0_18_RW0_wdata = RW0_wdata[151:144];
  assign mem_0_18_RW0_en = RW0_en;
  assign mem_0_18_RW0_wmode = RW0_wmode;
  assign mem_0_18_RW0_wmask = RW0_wmask[18];
  assign mem_0_19_RW0_addr = RW0_addr;
  assign mem_0_19_RW0_clk = RW0_clk;
  assign mem_0_19_RW0_wdata = RW0_wdata[159:152];
  assign mem_0_19_RW0_en = RW0_en;
  assign mem_0_19_RW0_wmode = RW0_wmode;
  assign mem_0_19_RW0_wmask = RW0_wmask[19];
  assign mem_0_20_RW0_addr = RW0_addr;
  assign mem_0_20_RW0_clk = RW0_clk;
  assign mem_0_20_RW0_wdata = RW0_wdata[167:160];
  assign mem_0_20_RW0_en = RW0_en;
  assign mem_0_20_RW0_wmode = RW0_wmode;
  assign mem_0_20_RW0_wmask = RW0_wmask[20];
  assign mem_0_21_RW0_addr = RW0_addr;
  assign mem_0_21_RW0_clk = RW0_clk;
  assign mem_0_21_RW0_wdata = RW0_wdata[175:168];
  assign mem_0_21_RW0_en = RW0_en;
  assign mem_0_21_RW0_wmode = RW0_wmode;
  assign mem_0_21_RW0_wmask = RW0_wmask[21];
  assign mem_0_22_RW0_addr = RW0_addr;
  assign mem_0_22_RW0_clk = RW0_clk;
  assign mem_0_22_RW0_wdata = RW0_wdata[183:176];
  assign mem_0_22_RW0_en = RW0_en;
  assign mem_0_22_RW0_wmode = RW0_wmode;
  assign mem_0_22_RW0_wmask = RW0_wmask[22];
  assign mem_0_23_RW0_addr = RW0_addr;
  assign mem_0_23_RW0_clk = RW0_clk;
  assign mem_0_23_RW0_wdata = RW0_wdata[191:184];
  assign mem_0_23_RW0_en = RW0_en;
  assign mem_0_23_RW0_wmode = RW0_wmode;
  assign mem_0_23_RW0_wmask = RW0_wmask[23];
  assign mem_0_24_RW0_addr = RW0_addr;
  assign mem_0_24_RW0_clk = RW0_clk;
  assign mem_0_24_RW0_wdata = RW0_wdata[199:192];
  assign mem_0_24_RW0_en = RW0_en;
  assign mem_0_24_RW0_wmode = RW0_wmode;
  assign mem_0_24_RW0_wmask = RW0_wmask[24];
  assign mem_0_25_RW0_addr = RW0_addr;
  assign mem_0_25_RW0_clk = RW0_clk;
  assign mem_0_25_RW0_wdata = RW0_wdata[207:200];
  assign mem_0_25_RW0_en = RW0_en;
  assign mem_0_25_RW0_wmode = RW0_wmode;
  assign mem_0_25_RW0_wmask = RW0_wmask[25];
  assign mem_0_26_RW0_addr = RW0_addr;
  assign mem_0_26_RW0_clk = RW0_clk;
  assign mem_0_26_RW0_wdata = RW0_wdata[215:208];
  assign mem_0_26_RW0_en = RW0_en;
  assign mem_0_26_RW0_wmode = RW0_wmode;
  assign mem_0_26_RW0_wmask = RW0_wmask[26];
  assign mem_0_27_RW0_addr = RW0_addr;
  assign mem_0_27_RW0_clk = RW0_clk;
  assign mem_0_27_RW0_wdata = RW0_wdata[223:216];
  assign mem_0_27_RW0_en = RW0_en;
  assign mem_0_27_RW0_wmode = RW0_wmode;
  assign mem_0_27_RW0_wmask = RW0_wmask[27];
  assign mem_0_28_RW0_addr = RW0_addr;
  assign mem_0_28_RW0_clk = RW0_clk;
  assign mem_0_28_RW0_wdata = RW0_wdata[231:224];
  assign mem_0_28_RW0_en = RW0_en;
  assign mem_0_28_RW0_wmode = RW0_wmode;
  assign mem_0_28_RW0_wmask = RW0_wmask[28];
  assign mem_0_29_RW0_addr = RW0_addr;
  assign mem_0_29_RW0_clk = RW0_clk;
  assign mem_0_29_RW0_wdata = RW0_wdata[239:232];
  assign mem_0_29_RW0_en = RW0_en;
  assign mem_0_29_RW0_wmode = RW0_wmode;
  assign mem_0_29_RW0_wmask = RW0_wmask[29];
  assign mem_0_30_RW0_addr = RW0_addr;
  assign mem_0_30_RW0_clk = RW0_clk;
  assign mem_0_30_RW0_wdata = RW0_wdata[247:240];
  assign mem_0_30_RW0_en = RW0_en;
  assign mem_0_30_RW0_wmode = RW0_wmode;
  assign mem_0_30_RW0_wmask = RW0_wmask[30];
  assign mem_0_31_RW0_addr = RW0_addr;
  assign mem_0_31_RW0_clk = RW0_clk;
  assign mem_0_31_RW0_wdata = RW0_wdata[255:248];
  assign mem_0_31_RW0_en = RW0_en;
  assign mem_0_31_RW0_wmode = RW0_wmode;
  assign mem_0_31_RW0_wmask = RW0_wmask[31];
endmodule
module tag_array_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [87:0] RW0_wdata,
  output [87:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input  [3:0]  RW0_wmask
);
  wire [5:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [21:0] mem_0_0_RW0_wdata;
  wire [21:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [5:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [21:0] mem_0_1_RW0_wdata;
  wire [21:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [5:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [21:0] mem_0_2_RW0_wdata;
  wire [21:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [5:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [21:0] mem_0_3_RW0_wdata;
  wire [21:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [21:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [21:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [21:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [21:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [43:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [65:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [87:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [43:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [65:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  split_tag_array_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[21:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[43:22];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[65:44];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[87:66];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
endmodule
module mem_ext(
  input  [11:0]  RW0_addr,
  input          RW0_clk,
  input  [127:0] RW0_wdata,
  output [127:0] RW0_rdata,
  input          RW0_en,
  input          RW0_wmode,
  input  [15:0]  RW0_wmask
);
  wire [11:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [7:0] mem_0_0_RW0_wdata;
  wire [7:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [11:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [7:0] mem_0_1_RW0_wdata;
  wire [7:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [11:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [7:0] mem_0_2_RW0_wdata;
  wire [7:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [11:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [7:0] mem_0_3_RW0_wdata;
  wire [7:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [11:0] mem_0_4_RW0_addr;
  wire  mem_0_4_RW0_clk;
  wire [7:0] mem_0_4_RW0_wdata;
  wire [7:0] mem_0_4_RW0_rdata;
  wire  mem_0_4_RW0_en;
  wire  mem_0_4_RW0_wmode;
  wire  mem_0_4_RW0_wmask;
  wire [11:0] mem_0_5_RW0_addr;
  wire  mem_0_5_RW0_clk;
  wire [7:0] mem_0_5_RW0_wdata;
  wire [7:0] mem_0_5_RW0_rdata;
  wire  mem_0_5_RW0_en;
  wire  mem_0_5_RW0_wmode;
  wire  mem_0_5_RW0_wmask;
  wire [11:0] mem_0_6_RW0_addr;
  wire  mem_0_6_RW0_clk;
  wire [7:0] mem_0_6_RW0_wdata;
  wire [7:0] mem_0_6_RW0_rdata;
  wire  mem_0_6_RW0_en;
  wire  mem_0_6_RW0_wmode;
  wire  mem_0_6_RW0_wmask;
  wire [11:0] mem_0_7_RW0_addr;
  wire  mem_0_7_RW0_clk;
  wire [7:0] mem_0_7_RW0_wdata;
  wire [7:0] mem_0_7_RW0_rdata;
  wire  mem_0_7_RW0_en;
  wire  mem_0_7_RW0_wmode;
  wire  mem_0_7_RW0_wmask;
  wire [11:0] mem_0_8_RW0_addr;
  wire  mem_0_8_RW0_clk;
  wire [7:0] mem_0_8_RW0_wdata;
  wire [7:0] mem_0_8_RW0_rdata;
  wire  mem_0_8_RW0_en;
  wire  mem_0_8_RW0_wmode;
  wire  mem_0_8_RW0_wmask;
  wire [11:0] mem_0_9_RW0_addr;
  wire  mem_0_9_RW0_clk;
  wire [7:0] mem_0_9_RW0_wdata;
  wire [7:0] mem_0_9_RW0_rdata;
  wire  mem_0_9_RW0_en;
  wire  mem_0_9_RW0_wmode;
  wire  mem_0_9_RW0_wmask;
  wire [11:0] mem_0_10_RW0_addr;
  wire  mem_0_10_RW0_clk;
  wire [7:0] mem_0_10_RW0_wdata;
  wire [7:0] mem_0_10_RW0_rdata;
  wire  mem_0_10_RW0_en;
  wire  mem_0_10_RW0_wmode;
  wire  mem_0_10_RW0_wmask;
  wire [11:0] mem_0_11_RW0_addr;
  wire  mem_0_11_RW0_clk;
  wire [7:0] mem_0_11_RW0_wdata;
  wire [7:0] mem_0_11_RW0_rdata;
  wire  mem_0_11_RW0_en;
  wire  mem_0_11_RW0_wmode;
  wire  mem_0_11_RW0_wmask;
  wire [11:0] mem_0_12_RW0_addr;
  wire  mem_0_12_RW0_clk;
  wire [7:0] mem_0_12_RW0_wdata;
  wire [7:0] mem_0_12_RW0_rdata;
  wire  mem_0_12_RW0_en;
  wire  mem_0_12_RW0_wmode;
  wire  mem_0_12_RW0_wmask;
  wire [11:0] mem_0_13_RW0_addr;
  wire  mem_0_13_RW0_clk;
  wire [7:0] mem_0_13_RW0_wdata;
  wire [7:0] mem_0_13_RW0_rdata;
  wire  mem_0_13_RW0_en;
  wire  mem_0_13_RW0_wmode;
  wire  mem_0_13_RW0_wmask;
  wire [11:0] mem_0_14_RW0_addr;
  wire  mem_0_14_RW0_clk;
  wire [7:0] mem_0_14_RW0_wdata;
  wire [7:0] mem_0_14_RW0_rdata;
  wire  mem_0_14_RW0_en;
  wire  mem_0_14_RW0_wmode;
  wire  mem_0_14_RW0_wmask;
  wire [11:0] mem_0_15_RW0_addr;
  wire  mem_0_15_RW0_clk;
  wire [7:0] mem_0_15_RW0_wdata;
  wire [7:0] mem_0_15_RW0_rdata;
  wire  mem_0_15_RW0_en;
  wire  mem_0_15_RW0_wmode;
  wire  mem_0_15_RW0_wmask;
  wire [7:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [7:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [7:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [7:0] RW0_rdata_0_4 = mem_0_4_RW0_rdata;
  wire [7:0] RW0_rdata_0_5 = mem_0_5_RW0_rdata;
  wire [7:0] RW0_rdata_0_6 = mem_0_6_RW0_rdata;
  wire [7:0] RW0_rdata_0_7 = mem_0_7_RW0_rdata;
  wire [7:0] RW0_rdata_0_8 = mem_0_8_RW0_rdata;
  wire [7:0] RW0_rdata_0_9 = mem_0_9_RW0_rdata;
  wire [7:0] RW0_rdata_0_10 = mem_0_10_RW0_rdata;
  wire [7:0] RW0_rdata_0_11 = mem_0_11_RW0_rdata;
  wire [7:0] RW0_rdata_0_12 = mem_0_12_RW0_rdata;
  wire [7:0] RW0_rdata_0_13 = mem_0_13_RW0_rdata;
  wire [7:0] RW0_rdata_0_14 = mem_0_14_RW0_rdata;
  wire [7:0] RW0_rdata_0_15 = mem_0_15_RW0_rdata;
  wire [15:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [31:0] _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [39:0] _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [47:0] _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [55:0] _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  wire [63:0] _GEN_6 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0};
  wire [71:0] _GEN_7 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,
    RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [79:0] _GEN_8 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,
    RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [87:0] _GEN_9 = {RW0_rdata_0_10,_GEN_8};
  wire [95:0] _GEN_10 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [103:0] _GEN_11 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [111:0] _GEN_12 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [119:0] _GEN_13 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [127:0] RW0_rdata_0 = {RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,
    _GEN_8};
  wire [15:0] _GEN_14 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_15 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [31:0] _GEN_16 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [39:0] _GEN_17 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [47:0] _GEN_18 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [55:0] _GEN_19 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0};
  wire [63:0] _GEN_20 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0};
  wire [71:0] _GEN_21 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,
    RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [79:0] _GEN_22 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,
    RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [87:0] _GEN_23 = {RW0_rdata_0_10,_GEN_8};
  wire [95:0] _GEN_24 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [103:0] _GEN_25 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [111:0] _GEN_26 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  wire [119:0] _GEN_27 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8};
  split_mem_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_mem_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_mem_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_mem_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_mem_ext mem_0_4 (
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_mem_ext mem_0_5 (
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_mem_ext mem_0_6 (
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_mem_ext mem_0_7 (
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  split_mem_ext mem_0_8 (
    .RW0_addr(mem_0_8_RW0_addr),
    .RW0_clk(mem_0_8_RW0_clk),
    .RW0_wdata(mem_0_8_RW0_wdata),
    .RW0_rdata(mem_0_8_RW0_rdata),
    .RW0_en(mem_0_8_RW0_en),
    .RW0_wmode(mem_0_8_RW0_wmode),
    .RW0_wmask(mem_0_8_RW0_wmask)
  );
  split_mem_ext mem_0_9 (
    .RW0_addr(mem_0_9_RW0_addr),
    .RW0_clk(mem_0_9_RW0_clk),
    .RW0_wdata(mem_0_9_RW0_wdata),
    .RW0_rdata(mem_0_9_RW0_rdata),
    .RW0_en(mem_0_9_RW0_en),
    .RW0_wmode(mem_0_9_RW0_wmode),
    .RW0_wmask(mem_0_9_RW0_wmask)
  );
  split_mem_ext mem_0_10 (
    .RW0_addr(mem_0_10_RW0_addr),
    .RW0_clk(mem_0_10_RW0_clk),
    .RW0_wdata(mem_0_10_RW0_wdata),
    .RW0_rdata(mem_0_10_RW0_rdata),
    .RW0_en(mem_0_10_RW0_en),
    .RW0_wmode(mem_0_10_RW0_wmode),
    .RW0_wmask(mem_0_10_RW0_wmask)
  );
  split_mem_ext mem_0_11 (
    .RW0_addr(mem_0_11_RW0_addr),
    .RW0_clk(mem_0_11_RW0_clk),
    .RW0_wdata(mem_0_11_RW0_wdata),
    .RW0_rdata(mem_0_11_RW0_rdata),
    .RW0_en(mem_0_11_RW0_en),
    .RW0_wmode(mem_0_11_RW0_wmode),
    .RW0_wmask(mem_0_11_RW0_wmask)
  );
  split_mem_ext mem_0_12 (
    .RW0_addr(mem_0_12_RW0_addr),
    .RW0_clk(mem_0_12_RW0_clk),
    .RW0_wdata(mem_0_12_RW0_wdata),
    .RW0_rdata(mem_0_12_RW0_rdata),
    .RW0_en(mem_0_12_RW0_en),
    .RW0_wmode(mem_0_12_RW0_wmode),
    .RW0_wmask(mem_0_12_RW0_wmask)
  );
  split_mem_ext mem_0_13 (
    .RW0_addr(mem_0_13_RW0_addr),
    .RW0_clk(mem_0_13_RW0_clk),
    .RW0_wdata(mem_0_13_RW0_wdata),
    .RW0_rdata(mem_0_13_RW0_rdata),
    .RW0_en(mem_0_13_RW0_en),
    .RW0_wmode(mem_0_13_RW0_wmode),
    .RW0_wmask(mem_0_13_RW0_wmask)
  );
  split_mem_ext mem_0_14 (
    .RW0_addr(mem_0_14_RW0_addr),
    .RW0_clk(mem_0_14_RW0_clk),
    .RW0_wdata(mem_0_14_RW0_wdata),
    .RW0_rdata(mem_0_14_RW0_rdata),
    .RW0_en(mem_0_14_RW0_en),
    .RW0_wmode(mem_0_14_RW0_wmode),
    .RW0_wmask(mem_0_14_RW0_wmask)
  );
  split_mem_ext mem_0_15 (
    .RW0_addr(mem_0_15_RW0_addr),
    .RW0_clk(mem_0_15_RW0_clk),
    .RW0_wdata(mem_0_15_RW0_wdata),
    .RW0_rdata(mem_0_15_RW0_rdata),
    .RW0_en(mem_0_15_RW0_en),
    .RW0_wmode(mem_0_15_RW0_wmode),
    .RW0_wmask(mem_0_15_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_15,_GEN_13};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[7:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[15:8];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[23:16];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[31:24];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
  assign mem_0_4_RW0_addr = RW0_addr;
  assign mem_0_4_RW0_clk = RW0_clk;
  assign mem_0_4_RW0_wdata = RW0_wdata[39:32];
  assign mem_0_4_RW0_en = RW0_en;
  assign mem_0_4_RW0_wmode = RW0_wmode;
  assign mem_0_4_RW0_wmask = RW0_wmask[4];
  assign mem_0_5_RW0_addr = RW0_addr;
  assign mem_0_5_RW0_clk = RW0_clk;
  assign mem_0_5_RW0_wdata = RW0_wdata[47:40];
  assign mem_0_5_RW0_en = RW0_en;
  assign mem_0_5_RW0_wmode = RW0_wmode;
  assign mem_0_5_RW0_wmask = RW0_wmask[5];
  assign mem_0_6_RW0_addr = RW0_addr;
  assign mem_0_6_RW0_clk = RW0_clk;
  assign mem_0_6_RW0_wdata = RW0_wdata[55:48];
  assign mem_0_6_RW0_en = RW0_en;
  assign mem_0_6_RW0_wmode = RW0_wmode;
  assign mem_0_6_RW0_wmask = RW0_wmask[6];
  assign mem_0_7_RW0_addr = RW0_addr;
  assign mem_0_7_RW0_clk = RW0_clk;
  assign mem_0_7_RW0_wdata = RW0_wdata[63:56];
  assign mem_0_7_RW0_en = RW0_en;
  assign mem_0_7_RW0_wmode = RW0_wmode;
  assign mem_0_7_RW0_wmask = RW0_wmask[7];
  assign mem_0_8_RW0_addr = RW0_addr;
  assign mem_0_8_RW0_clk = RW0_clk;
  assign mem_0_8_RW0_wdata = RW0_wdata[71:64];
  assign mem_0_8_RW0_en = RW0_en;
  assign mem_0_8_RW0_wmode = RW0_wmode;
  assign mem_0_8_RW0_wmask = RW0_wmask[8];
  assign mem_0_9_RW0_addr = RW0_addr;
  assign mem_0_9_RW0_clk = RW0_clk;
  assign mem_0_9_RW0_wdata = RW0_wdata[79:72];
  assign mem_0_9_RW0_en = RW0_en;
  assign mem_0_9_RW0_wmode = RW0_wmode;
  assign mem_0_9_RW0_wmask = RW0_wmask[9];
  assign mem_0_10_RW0_addr = RW0_addr;
  assign mem_0_10_RW0_clk = RW0_clk;
  assign mem_0_10_RW0_wdata = RW0_wdata[87:80];
  assign mem_0_10_RW0_en = RW0_en;
  assign mem_0_10_RW0_wmode = RW0_wmode;
  assign mem_0_10_RW0_wmask = RW0_wmask[10];
  assign mem_0_11_RW0_addr = RW0_addr;
  assign mem_0_11_RW0_clk = RW0_clk;
  assign mem_0_11_RW0_wdata = RW0_wdata[95:88];
  assign mem_0_11_RW0_en = RW0_en;
  assign mem_0_11_RW0_wmode = RW0_wmode;
  assign mem_0_11_RW0_wmask = RW0_wmask[11];
  assign mem_0_12_RW0_addr = RW0_addr;
  assign mem_0_12_RW0_clk = RW0_clk;
  assign mem_0_12_RW0_wdata = RW0_wdata[103:96];
  assign mem_0_12_RW0_en = RW0_en;
  assign mem_0_12_RW0_wmode = RW0_wmode;
  assign mem_0_12_RW0_wmask = RW0_wmask[12];
  assign mem_0_13_RW0_addr = RW0_addr;
  assign mem_0_13_RW0_clk = RW0_clk;
  assign mem_0_13_RW0_wdata = RW0_wdata[111:104];
  assign mem_0_13_RW0_en = RW0_en;
  assign mem_0_13_RW0_wmode = RW0_wmode;
  assign mem_0_13_RW0_wmask = RW0_wmask[13];
  assign mem_0_14_RW0_addr = RW0_addr;
  assign mem_0_14_RW0_clk = RW0_clk;
  assign mem_0_14_RW0_wdata = RW0_wdata[119:112];
  assign mem_0_14_RW0_en = RW0_en;
  assign mem_0_14_RW0_wmode = RW0_wmode;
  assign mem_0_14_RW0_wmask = RW0_wmask[14];
  assign mem_0_15_RW0_addr = RW0_addr;
  assign mem_0_15_RW0_clk = RW0_clk;
  assign mem_0_15_RW0_wdata = RW0_wdata[127:120];
  assign mem_0_15_RW0_en = RW0_en;
  assign mem_0_15_RW0_wmode = RW0_wmode;
  assign mem_0_15_RW0_wmask = RW0_wmask[15];
endmodule
module mem_0_ext(
  input  [8:0]   R0_addr,
  input          R0_clk,
  output [511:0] R0_data,
  input          R0_en,
  input  [8:0]   W0_addr,
  input          W0_clk,
  input  [511:0] W0_data,
  input          W0_en,
  input  [63:0]  W0_mask
);
  wire [8:0] mem_0_0_R0_addr;
  wire  mem_0_0_R0_clk;
  wire [7:0] mem_0_0_R0_data;
  wire  mem_0_0_R0_en;
  wire [8:0] mem_0_0_W0_addr;
  wire  mem_0_0_W0_clk;
  wire [7:0] mem_0_0_W0_data;
  wire  mem_0_0_W0_en;
  wire  mem_0_0_W0_mask;
  wire [8:0] mem_0_1_R0_addr;
  wire  mem_0_1_R0_clk;
  wire [7:0] mem_0_1_R0_data;
  wire  mem_0_1_R0_en;
  wire [8:0] mem_0_1_W0_addr;
  wire  mem_0_1_W0_clk;
  wire [7:0] mem_0_1_W0_data;
  wire  mem_0_1_W0_en;
  wire  mem_0_1_W0_mask;
  wire [8:0] mem_0_2_R0_addr;
  wire  mem_0_2_R0_clk;
  wire [7:0] mem_0_2_R0_data;
  wire  mem_0_2_R0_en;
  wire [8:0] mem_0_2_W0_addr;
  wire  mem_0_2_W0_clk;
  wire [7:0] mem_0_2_W0_data;
  wire  mem_0_2_W0_en;
  wire  mem_0_2_W0_mask;
  wire [8:0] mem_0_3_R0_addr;
  wire  mem_0_3_R0_clk;
  wire [7:0] mem_0_3_R0_data;
  wire  mem_0_3_R0_en;
  wire [8:0] mem_0_3_W0_addr;
  wire  mem_0_3_W0_clk;
  wire [7:0] mem_0_3_W0_data;
  wire  mem_0_3_W0_en;
  wire  mem_0_3_W0_mask;
  wire [8:0] mem_0_4_R0_addr;
  wire  mem_0_4_R0_clk;
  wire [7:0] mem_0_4_R0_data;
  wire  mem_0_4_R0_en;
  wire [8:0] mem_0_4_W0_addr;
  wire  mem_0_4_W0_clk;
  wire [7:0] mem_0_4_W0_data;
  wire  mem_0_4_W0_en;
  wire  mem_0_4_W0_mask;
  wire [8:0] mem_0_5_R0_addr;
  wire  mem_0_5_R0_clk;
  wire [7:0] mem_0_5_R0_data;
  wire  mem_0_5_R0_en;
  wire [8:0] mem_0_5_W0_addr;
  wire  mem_0_5_W0_clk;
  wire [7:0] mem_0_5_W0_data;
  wire  mem_0_5_W0_en;
  wire  mem_0_5_W0_mask;
  wire [8:0] mem_0_6_R0_addr;
  wire  mem_0_6_R0_clk;
  wire [7:0] mem_0_6_R0_data;
  wire  mem_0_6_R0_en;
  wire [8:0] mem_0_6_W0_addr;
  wire  mem_0_6_W0_clk;
  wire [7:0] mem_0_6_W0_data;
  wire  mem_0_6_W0_en;
  wire  mem_0_6_W0_mask;
  wire [8:0] mem_0_7_R0_addr;
  wire  mem_0_7_R0_clk;
  wire [7:0] mem_0_7_R0_data;
  wire  mem_0_7_R0_en;
  wire [8:0] mem_0_7_W0_addr;
  wire  mem_0_7_W0_clk;
  wire [7:0] mem_0_7_W0_data;
  wire  mem_0_7_W0_en;
  wire  mem_0_7_W0_mask;
  wire [8:0] mem_0_8_R0_addr;
  wire  mem_0_8_R0_clk;
  wire [7:0] mem_0_8_R0_data;
  wire  mem_0_8_R0_en;
  wire [8:0] mem_0_8_W0_addr;
  wire  mem_0_8_W0_clk;
  wire [7:0] mem_0_8_W0_data;
  wire  mem_0_8_W0_en;
  wire  mem_0_8_W0_mask;
  wire [8:0] mem_0_9_R0_addr;
  wire  mem_0_9_R0_clk;
  wire [7:0] mem_0_9_R0_data;
  wire  mem_0_9_R0_en;
  wire [8:0] mem_0_9_W0_addr;
  wire  mem_0_9_W0_clk;
  wire [7:0] mem_0_9_W0_data;
  wire  mem_0_9_W0_en;
  wire  mem_0_9_W0_mask;
  wire [8:0] mem_0_10_R0_addr;
  wire  mem_0_10_R0_clk;
  wire [7:0] mem_0_10_R0_data;
  wire  mem_0_10_R0_en;
  wire [8:0] mem_0_10_W0_addr;
  wire  mem_0_10_W0_clk;
  wire [7:0] mem_0_10_W0_data;
  wire  mem_0_10_W0_en;
  wire  mem_0_10_W0_mask;
  wire [8:0] mem_0_11_R0_addr;
  wire  mem_0_11_R0_clk;
  wire [7:0] mem_0_11_R0_data;
  wire  mem_0_11_R0_en;
  wire [8:0] mem_0_11_W0_addr;
  wire  mem_0_11_W0_clk;
  wire [7:0] mem_0_11_W0_data;
  wire  mem_0_11_W0_en;
  wire  mem_0_11_W0_mask;
  wire [8:0] mem_0_12_R0_addr;
  wire  mem_0_12_R0_clk;
  wire [7:0] mem_0_12_R0_data;
  wire  mem_0_12_R0_en;
  wire [8:0] mem_0_12_W0_addr;
  wire  mem_0_12_W0_clk;
  wire [7:0] mem_0_12_W0_data;
  wire  mem_0_12_W0_en;
  wire  mem_0_12_W0_mask;
  wire [8:0] mem_0_13_R0_addr;
  wire  mem_0_13_R0_clk;
  wire [7:0] mem_0_13_R0_data;
  wire  mem_0_13_R0_en;
  wire [8:0] mem_0_13_W0_addr;
  wire  mem_0_13_W0_clk;
  wire [7:0] mem_0_13_W0_data;
  wire  mem_0_13_W0_en;
  wire  mem_0_13_W0_mask;
  wire [8:0] mem_0_14_R0_addr;
  wire  mem_0_14_R0_clk;
  wire [7:0] mem_0_14_R0_data;
  wire  mem_0_14_R0_en;
  wire [8:0] mem_0_14_W0_addr;
  wire  mem_0_14_W0_clk;
  wire [7:0] mem_0_14_W0_data;
  wire  mem_0_14_W0_en;
  wire  mem_0_14_W0_mask;
  wire [8:0] mem_0_15_R0_addr;
  wire  mem_0_15_R0_clk;
  wire [7:0] mem_0_15_R0_data;
  wire  mem_0_15_R0_en;
  wire [8:0] mem_0_15_W0_addr;
  wire  mem_0_15_W0_clk;
  wire [7:0] mem_0_15_W0_data;
  wire  mem_0_15_W0_en;
  wire  mem_0_15_W0_mask;
  wire [8:0] mem_0_16_R0_addr;
  wire  mem_0_16_R0_clk;
  wire [7:0] mem_0_16_R0_data;
  wire  mem_0_16_R0_en;
  wire [8:0] mem_0_16_W0_addr;
  wire  mem_0_16_W0_clk;
  wire [7:0] mem_0_16_W0_data;
  wire  mem_0_16_W0_en;
  wire  mem_0_16_W0_mask;
  wire [8:0] mem_0_17_R0_addr;
  wire  mem_0_17_R0_clk;
  wire [7:0] mem_0_17_R0_data;
  wire  mem_0_17_R0_en;
  wire [8:0] mem_0_17_W0_addr;
  wire  mem_0_17_W0_clk;
  wire [7:0] mem_0_17_W0_data;
  wire  mem_0_17_W0_en;
  wire  mem_0_17_W0_mask;
  wire [8:0] mem_0_18_R0_addr;
  wire  mem_0_18_R0_clk;
  wire [7:0] mem_0_18_R0_data;
  wire  mem_0_18_R0_en;
  wire [8:0] mem_0_18_W0_addr;
  wire  mem_0_18_W0_clk;
  wire [7:0] mem_0_18_W0_data;
  wire  mem_0_18_W0_en;
  wire  mem_0_18_W0_mask;
  wire [8:0] mem_0_19_R0_addr;
  wire  mem_0_19_R0_clk;
  wire [7:0] mem_0_19_R0_data;
  wire  mem_0_19_R0_en;
  wire [8:0] mem_0_19_W0_addr;
  wire  mem_0_19_W0_clk;
  wire [7:0] mem_0_19_W0_data;
  wire  mem_0_19_W0_en;
  wire  mem_0_19_W0_mask;
  wire [8:0] mem_0_20_R0_addr;
  wire  mem_0_20_R0_clk;
  wire [7:0] mem_0_20_R0_data;
  wire  mem_0_20_R0_en;
  wire [8:0] mem_0_20_W0_addr;
  wire  mem_0_20_W0_clk;
  wire [7:0] mem_0_20_W0_data;
  wire  mem_0_20_W0_en;
  wire  mem_0_20_W0_mask;
  wire [8:0] mem_0_21_R0_addr;
  wire  mem_0_21_R0_clk;
  wire [7:0] mem_0_21_R0_data;
  wire  mem_0_21_R0_en;
  wire [8:0] mem_0_21_W0_addr;
  wire  mem_0_21_W0_clk;
  wire [7:0] mem_0_21_W0_data;
  wire  mem_0_21_W0_en;
  wire  mem_0_21_W0_mask;
  wire [8:0] mem_0_22_R0_addr;
  wire  mem_0_22_R0_clk;
  wire [7:0] mem_0_22_R0_data;
  wire  mem_0_22_R0_en;
  wire [8:0] mem_0_22_W0_addr;
  wire  mem_0_22_W0_clk;
  wire [7:0] mem_0_22_W0_data;
  wire  mem_0_22_W0_en;
  wire  mem_0_22_W0_mask;
  wire [8:0] mem_0_23_R0_addr;
  wire  mem_0_23_R0_clk;
  wire [7:0] mem_0_23_R0_data;
  wire  mem_0_23_R0_en;
  wire [8:0] mem_0_23_W0_addr;
  wire  mem_0_23_W0_clk;
  wire [7:0] mem_0_23_W0_data;
  wire  mem_0_23_W0_en;
  wire  mem_0_23_W0_mask;
  wire [8:0] mem_0_24_R0_addr;
  wire  mem_0_24_R0_clk;
  wire [7:0] mem_0_24_R0_data;
  wire  mem_0_24_R0_en;
  wire [8:0] mem_0_24_W0_addr;
  wire  mem_0_24_W0_clk;
  wire [7:0] mem_0_24_W0_data;
  wire  mem_0_24_W0_en;
  wire  mem_0_24_W0_mask;
  wire [8:0] mem_0_25_R0_addr;
  wire  mem_0_25_R0_clk;
  wire [7:0] mem_0_25_R0_data;
  wire  mem_0_25_R0_en;
  wire [8:0] mem_0_25_W0_addr;
  wire  mem_0_25_W0_clk;
  wire [7:0] mem_0_25_W0_data;
  wire  mem_0_25_W0_en;
  wire  mem_0_25_W0_mask;
  wire [8:0] mem_0_26_R0_addr;
  wire  mem_0_26_R0_clk;
  wire [7:0] mem_0_26_R0_data;
  wire  mem_0_26_R0_en;
  wire [8:0] mem_0_26_W0_addr;
  wire  mem_0_26_W0_clk;
  wire [7:0] mem_0_26_W0_data;
  wire  mem_0_26_W0_en;
  wire  mem_0_26_W0_mask;
  wire [8:0] mem_0_27_R0_addr;
  wire  mem_0_27_R0_clk;
  wire [7:0] mem_0_27_R0_data;
  wire  mem_0_27_R0_en;
  wire [8:0] mem_0_27_W0_addr;
  wire  mem_0_27_W0_clk;
  wire [7:0] mem_0_27_W0_data;
  wire  mem_0_27_W0_en;
  wire  mem_0_27_W0_mask;
  wire [8:0] mem_0_28_R0_addr;
  wire  mem_0_28_R0_clk;
  wire [7:0] mem_0_28_R0_data;
  wire  mem_0_28_R0_en;
  wire [8:0] mem_0_28_W0_addr;
  wire  mem_0_28_W0_clk;
  wire [7:0] mem_0_28_W0_data;
  wire  mem_0_28_W0_en;
  wire  mem_0_28_W0_mask;
  wire [8:0] mem_0_29_R0_addr;
  wire  mem_0_29_R0_clk;
  wire [7:0] mem_0_29_R0_data;
  wire  mem_0_29_R0_en;
  wire [8:0] mem_0_29_W0_addr;
  wire  mem_0_29_W0_clk;
  wire [7:0] mem_0_29_W0_data;
  wire  mem_0_29_W0_en;
  wire  mem_0_29_W0_mask;
  wire [8:0] mem_0_30_R0_addr;
  wire  mem_0_30_R0_clk;
  wire [7:0] mem_0_30_R0_data;
  wire  mem_0_30_R0_en;
  wire [8:0] mem_0_30_W0_addr;
  wire  mem_0_30_W0_clk;
  wire [7:0] mem_0_30_W0_data;
  wire  mem_0_30_W0_en;
  wire  mem_0_30_W0_mask;
  wire [8:0] mem_0_31_R0_addr;
  wire  mem_0_31_R0_clk;
  wire [7:0] mem_0_31_R0_data;
  wire  mem_0_31_R0_en;
  wire [8:0] mem_0_31_W0_addr;
  wire  mem_0_31_W0_clk;
  wire [7:0] mem_0_31_W0_data;
  wire  mem_0_31_W0_en;
  wire  mem_0_31_W0_mask;
  wire [8:0] mem_0_32_R0_addr;
  wire  mem_0_32_R0_clk;
  wire [7:0] mem_0_32_R0_data;
  wire  mem_0_32_R0_en;
  wire [8:0] mem_0_32_W0_addr;
  wire  mem_0_32_W0_clk;
  wire [7:0] mem_0_32_W0_data;
  wire  mem_0_32_W0_en;
  wire  mem_0_32_W0_mask;
  wire [8:0] mem_0_33_R0_addr;
  wire  mem_0_33_R0_clk;
  wire [7:0] mem_0_33_R0_data;
  wire  mem_0_33_R0_en;
  wire [8:0] mem_0_33_W0_addr;
  wire  mem_0_33_W0_clk;
  wire [7:0] mem_0_33_W0_data;
  wire  mem_0_33_W0_en;
  wire  mem_0_33_W0_mask;
  wire [8:0] mem_0_34_R0_addr;
  wire  mem_0_34_R0_clk;
  wire [7:0] mem_0_34_R0_data;
  wire  mem_0_34_R0_en;
  wire [8:0] mem_0_34_W0_addr;
  wire  mem_0_34_W0_clk;
  wire [7:0] mem_0_34_W0_data;
  wire  mem_0_34_W0_en;
  wire  mem_0_34_W0_mask;
  wire [8:0] mem_0_35_R0_addr;
  wire  mem_0_35_R0_clk;
  wire [7:0] mem_0_35_R0_data;
  wire  mem_0_35_R0_en;
  wire [8:0] mem_0_35_W0_addr;
  wire  mem_0_35_W0_clk;
  wire [7:0] mem_0_35_W0_data;
  wire  mem_0_35_W0_en;
  wire  mem_0_35_W0_mask;
  wire [8:0] mem_0_36_R0_addr;
  wire  mem_0_36_R0_clk;
  wire [7:0] mem_0_36_R0_data;
  wire  mem_0_36_R0_en;
  wire [8:0] mem_0_36_W0_addr;
  wire  mem_0_36_W0_clk;
  wire [7:0] mem_0_36_W0_data;
  wire  mem_0_36_W0_en;
  wire  mem_0_36_W0_mask;
  wire [8:0] mem_0_37_R0_addr;
  wire  mem_0_37_R0_clk;
  wire [7:0] mem_0_37_R0_data;
  wire  mem_0_37_R0_en;
  wire [8:0] mem_0_37_W0_addr;
  wire  mem_0_37_W0_clk;
  wire [7:0] mem_0_37_W0_data;
  wire  mem_0_37_W0_en;
  wire  mem_0_37_W0_mask;
  wire [8:0] mem_0_38_R0_addr;
  wire  mem_0_38_R0_clk;
  wire [7:0] mem_0_38_R0_data;
  wire  mem_0_38_R0_en;
  wire [8:0] mem_0_38_W0_addr;
  wire  mem_0_38_W0_clk;
  wire [7:0] mem_0_38_W0_data;
  wire  mem_0_38_W0_en;
  wire  mem_0_38_W0_mask;
  wire [8:0] mem_0_39_R0_addr;
  wire  mem_0_39_R0_clk;
  wire [7:0] mem_0_39_R0_data;
  wire  mem_0_39_R0_en;
  wire [8:0] mem_0_39_W0_addr;
  wire  mem_0_39_W0_clk;
  wire [7:0] mem_0_39_W0_data;
  wire  mem_0_39_W0_en;
  wire  mem_0_39_W0_mask;
  wire [8:0] mem_0_40_R0_addr;
  wire  mem_0_40_R0_clk;
  wire [7:0] mem_0_40_R0_data;
  wire  mem_0_40_R0_en;
  wire [8:0] mem_0_40_W0_addr;
  wire  mem_0_40_W0_clk;
  wire [7:0] mem_0_40_W0_data;
  wire  mem_0_40_W0_en;
  wire  mem_0_40_W0_mask;
  wire [8:0] mem_0_41_R0_addr;
  wire  mem_0_41_R0_clk;
  wire [7:0] mem_0_41_R0_data;
  wire  mem_0_41_R0_en;
  wire [8:0] mem_0_41_W0_addr;
  wire  mem_0_41_W0_clk;
  wire [7:0] mem_0_41_W0_data;
  wire  mem_0_41_W0_en;
  wire  mem_0_41_W0_mask;
  wire [8:0] mem_0_42_R0_addr;
  wire  mem_0_42_R0_clk;
  wire [7:0] mem_0_42_R0_data;
  wire  mem_0_42_R0_en;
  wire [8:0] mem_0_42_W0_addr;
  wire  mem_0_42_W0_clk;
  wire [7:0] mem_0_42_W0_data;
  wire  mem_0_42_W0_en;
  wire  mem_0_42_W0_mask;
  wire [8:0] mem_0_43_R0_addr;
  wire  mem_0_43_R0_clk;
  wire [7:0] mem_0_43_R0_data;
  wire  mem_0_43_R0_en;
  wire [8:0] mem_0_43_W0_addr;
  wire  mem_0_43_W0_clk;
  wire [7:0] mem_0_43_W0_data;
  wire  mem_0_43_W0_en;
  wire  mem_0_43_W0_mask;
  wire [8:0] mem_0_44_R0_addr;
  wire  mem_0_44_R0_clk;
  wire [7:0] mem_0_44_R0_data;
  wire  mem_0_44_R0_en;
  wire [8:0] mem_0_44_W0_addr;
  wire  mem_0_44_W0_clk;
  wire [7:0] mem_0_44_W0_data;
  wire  mem_0_44_W0_en;
  wire  mem_0_44_W0_mask;
  wire [8:0] mem_0_45_R0_addr;
  wire  mem_0_45_R0_clk;
  wire [7:0] mem_0_45_R0_data;
  wire  mem_0_45_R0_en;
  wire [8:0] mem_0_45_W0_addr;
  wire  mem_0_45_W0_clk;
  wire [7:0] mem_0_45_W0_data;
  wire  mem_0_45_W0_en;
  wire  mem_0_45_W0_mask;
  wire [8:0] mem_0_46_R0_addr;
  wire  mem_0_46_R0_clk;
  wire [7:0] mem_0_46_R0_data;
  wire  mem_0_46_R0_en;
  wire [8:0] mem_0_46_W0_addr;
  wire  mem_0_46_W0_clk;
  wire [7:0] mem_0_46_W0_data;
  wire  mem_0_46_W0_en;
  wire  mem_0_46_W0_mask;
  wire [8:0] mem_0_47_R0_addr;
  wire  mem_0_47_R0_clk;
  wire [7:0] mem_0_47_R0_data;
  wire  mem_0_47_R0_en;
  wire [8:0] mem_0_47_W0_addr;
  wire  mem_0_47_W0_clk;
  wire [7:0] mem_0_47_W0_data;
  wire  mem_0_47_W0_en;
  wire  mem_0_47_W0_mask;
  wire [8:0] mem_0_48_R0_addr;
  wire  mem_0_48_R0_clk;
  wire [7:0] mem_0_48_R0_data;
  wire  mem_0_48_R0_en;
  wire [8:0] mem_0_48_W0_addr;
  wire  mem_0_48_W0_clk;
  wire [7:0] mem_0_48_W0_data;
  wire  mem_0_48_W0_en;
  wire  mem_0_48_W0_mask;
  wire [8:0] mem_0_49_R0_addr;
  wire  mem_0_49_R0_clk;
  wire [7:0] mem_0_49_R0_data;
  wire  mem_0_49_R0_en;
  wire [8:0] mem_0_49_W0_addr;
  wire  mem_0_49_W0_clk;
  wire [7:0] mem_0_49_W0_data;
  wire  mem_0_49_W0_en;
  wire  mem_0_49_W0_mask;
  wire [8:0] mem_0_50_R0_addr;
  wire  mem_0_50_R0_clk;
  wire [7:0] mem_0_50_R0_data;
  wire  mem_0_50_R0_en;
  wire [8:0] mem_0_50_W0_addr;
  wire  mem_0_50_W0_clk;
  wire [7:0] mem_0_50_W0_data;
  wire  mem_0_50_W0_en;
  wire  mem_0_50_W0_mask;
  wire [8:0] mem_0_51_R0_addr;
  wire  mem_0_51_R0_clk;
  wire [7:0] mem_0_51_R0_data;
  wire  mem_0_51_R0_en;
  wire [8:0] mem_0_51_W0_addr;
  wire  mem_0_51_W0_clk;
  wire [7:0] mem_0_51_W0_data;
  wire  mem_0_51_W0_en;
  wire  mem_0_51_W0_mask;
  wire [8:0] mem_0_52_R0_addr;
  wire  mem_0_52_R0_clk;
  wire [7:0] mem_0_52_R0_data;
  wire  mem_0_52_R0_en;
  wire [8:0] mem_0_52_W0_addr;
  wire  mem_0_52_W0_clk;
  wire [7:0] mem_0_52_W0_data;
  wire  mem_0_52_W0_en;
  wire  mem_0_52_W0_mask;
  wire [8:0] mem_0_53_R0_addr;
  wire  mem_0_53_R0_clk;
  wire [7:0] mem_0_53_R0_data;
  wire  mem_0_53_R0_en;
  wire [8:0] mem_0_53_W0_addr;
  wire  mem_0_53_W0_clk;
  wire [7:0] mem_0_53_W0_data;
  wire  mem_0_53_W0_en;
  wire  mem_0_53_W0_mask;
  wire [8:0] mem_0_54_R0_addr;
  wire  mem_0_54_R0_clk;
  wire [7:0] mem_0_54_R0_data;
  wire  mem_0_54_R0_en;
  wire [8:0] mem_0_54_W0_addr;
  wire  mem_0_54_W0_clk;
  wire [7:0] mem_0_54_W0_data;
  wire  mem_0_54_W0_en;
  wire  mem_0_54_W0_mask;
  wire [8:0] mem_0_55_R0_addr;
  wire  mem_0_55_R0_clk;
  wire [7:0] mem_0_55_R0_data;
  wire  mem_0_55_R0_en;
  wire [8:0] mem_0_55_W0_addr;
  wire  mem_0_55_W0_clk;
  wire [7:0] mem_0_55_W0_data;
  wire  mem_0_55_W0_en;
  wire  mem_0_55_W0_mask;
  wire [8:0] mem_0_56_R0_addr;
  wire  mem_0_56_R0_clk;
  wire [7:0] mem_0_56_R0_data;
  wire  mem_0_56_R0_en;
  wire [8:0] mem_0_56_W0_addr;
  wire  mem_0_56_W0_clk;
  wire [7:0] mem_0_56_W0_data;
  wire  mem_0_56_W0_en;
  wire  mem_0_56_W0_mask;
  wire [8:0] mem_0_57_R0_addr;
  wire  mem_0_57_R0_clk;
  wire [7:0] mem_0_57_R0_data;
  wire  mem_0_57_R0_en;
  wire [8:0] mem_0_57_W0_addr;
  wire  mem_0_57_W0_clk;
  wire [7:0] mem_0_57_W0_data;
  wire  mem_0_57_W0_en;
  wire  mem_0_57_W0_mask;
  wire [8:0] mem_0_58_R0_addr;
  wire  mem_0_58_R0_clk;
  wire [7:0] mem_0_58_R0_data;
  wire  mem_0_58_R0_en;
  wire [8:0] mem_0_58_W0_addr;
  wire  mem_0_58_W0_clk;
  wire [7:0] mem_0_58_W0_data;
  wire  mem_0_58_W0_en;
  wire  mem_0_58_W0_mask;
  wire [8:0] mem_0_59_R0_addr;
  wire  mem_0_59_R0_clk;
  wire [7:0] mem_0_59_R0_data;
  wire  mem_0_59_R0_en;
  wire [8:0] mem_0_59_W0_addr;
  wire  mem_0_59_W0_clk;
  wire [7:0] mem_0_59_W0_data;
  wire  mem_0_59_W0_en;
  wire  mem_0_59_W0_mask;
  wire [8:0] mem_0_60_R0_addr;
  wire  mem_0_60_R0_clk;
  wire [7:0] mem_0_60_R0_data;
  wire  mem_0_60_R0_en;
  wire [8:0] mem_0_60_W0_addr;
  wire  mem_0_60_W0_clk;
  wire [7:0] mem_0_60_W0_data;
  wire  mem_0_60_W0_en;
  wire  mem_0_60_W0_mask;
  wire [8:0] mem_0_61_R0_addr;
  wire  mem_0_61_R0_clk;
  wire [7:0] mem_0_61_R0_data;
  wire  mem_0_61_R0_en;
  wire [8:0] mem_0_61_W0_addr;
  wire  mem_0_61_W0_clk;
  wire [7:0] mem_0_61_W0_data;
  wire  mem_0_61_W0_en;
  wire  mem_0_61_W0_mask;
  wire [8:0] mem_0_62_R0_addr;
  wire  mem_0_62_R0_clk;
  wire [7:0] mem_0_62_R0_data;
  wire  mem_0_62_R0_en;
  wire [8:0] mem_0_62_W0_addr;
  wire  mem_0_62_W0_clk;
  wire [7:0] mem_0_62_W0_data;
  wire  mem_0_62_W0_en;
  wire  mem_0_62_W0_mask;
  wire [8:0] mem_0_63_R0_addr;
  wire  mem_0_63_R0_clk;
  wire [7:0] mem_0_63_R0_data;
  wire  mem_0_63_R0_en;
  wire [8:0] mem_0_63_W0_addr;
  wire  mem_0_63_W0_clk;
  wire [7:0] mem_0_63_W0_data;
  wire  mem_0_63_W0_en;
  wire  mem_0_63_W0_mask;
  wire [7:0] R0_data_0_0 = mem_0_0_R0_data;
  wire [7:0] R0_data_0_1 = mem_0_1_R0_data;
  wire [7:0] R0_data_0_2 = mem_0_2_R0_data;
  wire [7:0] R0_data_0_3 = mem_0_3_R0_data;
  wire [7:0] R0_data_0_4 = mem_0_4_R0_data;
  wire [7:0] R0_data_0_5 = mem_0_5_R0_data;
  wire [7:0] R0_data_0_6 = mem_0_6_R0_data;
  wire [7:0] R0_data_0_7 = mem_0_7_R0_data;
  wire [7:0] R0_data_0_8 = mem_0_8_R0_data;
  wire [7:0] R0_data_0_9 = mem_0_9_R0_data;
  wire [7:0] R0_data_0_10 = mem_0_10_R0_data;
  wire [7:0] R0_data_0_11 = mem_0_11_R0_data;
  wire [7:0] R0_data_0_12 = mem_0_12_R0_data;
  wire [7:0] R0_data_0_13 = mem_0_13_R0_data;
  wire [7:0] R0_data_0_14 = mem_0_14_R0_data;
  wire [7:0] R0_data_0_15 = mem_0_15_R0_data;
  wire [7:0] R0_data_0_16 = mem_0_16_R0_data;
  wire [7:0] R0_data_0_17 = mem_0_17_R0_data;
  wire [7:0] R0_data_0_18 = mem_0_18_R0_data;
  wire [7:0] R0_data_0_19 = mem_0_19_R0_data;
  wire [7:0] R0_data_0_20 = mem_0_20_R0_data;
  wire [7:0] R0_data_0_21 = mem_0_21_R0_data;
  wire [7:0] R0_data_0_22 = mem_0_22_R0_data;
  wire [7:0] R0_data_0_23 = mem_0_23_R0_data;
  wire [7:0] R0_data_0_24 = mem_0_24_R0_data;
  wire [7:0] R0_data_0_25 = mem_0_25_R0_data;
  wire [7:0] R0_data_0_26 = mem_0_26_R0_data;
  wire [7:0] R0_data_0_27 = mem_0_27_R0_data;
  wire [7:0] R0_data_0_28 = mem_0_28_R0_data;
  wire [7:0] R0_data_0_29 = mem_0_29_R0_data;
  wire [7:0] R0_data_0_30 = mem_0_30_R0_data;
  wire [7:0] R0_data_0_31 = mem_0_31_R0_data;
  wire [7:0] R0_data_0_32 = mem_0_32_R0_data;
  wire [7:0] R0_data_0_33 = mem_0_33_R0_data;
  wire [7:0] R0_data_0_34 = mem_0_34_R0_data;
  wire [7:0] R0_data_0_35 = mem_0_35_R0_data;
  wire [7:0] R0_data_0_36 = mem_0_36_R0_data;
  wire [7:0] R0_data_0_37 = mem_0_37_R0_data;
  wire [7:0] R0_data_0_38 = mem_0_38_R0_data;
  wire [7:0] R0_data_0_39 = mem_0_39_R0_data;
  wire [7:0] R0_data_0_40 = mem_0_40_R0_data;
  wire [7:0] R0_data_0_41 = mem_0_41_R0_data;
  wire [7:0] R0_data_0_42 = mem_0_42_R0_data;
  wire [7:0] R0_data_0_43 = mem_0_43_R0_data;
  wire [7:0] R0_data_0_44 = mem_0_44_R0_data;
  wire [7:0] R0_data_0_45 = mem_0_45_R0_data;
  wire [7:0] R0_data_0_46 = mem_0_46_R0_data;
  wire [7:0] R0_data_0_47 = mem_0_47_R0_data;
  wire [7:0] R0_data_0_48 = mem_0_48_R0_data;
  wire [7:0] R0_data_0_49 = mem_0_49_R0_data;
  wire [7:0] R0_data_0_50 = mem_0_50_R0_data;
  wire [7:0] R0_data_0_51 = mem_0_51_R0_data;
  wire [7:0] R0_data_0_52 = mem_0_52_R0_data;
  wire [7:0] R0_data_0_53 = mem_0_53_R0_data;
  wire [7:0] R0_data_0_54 = mem_0_54_R0_data;
  wire [7:0] R0_data_0_55 = mem_0_55_R0_data;
  wire [7:0] R0_data_0_56 = mem_0_56_R0_data;
  wire [7:0] R0_data_0_57 = mem_0_57_R0_data;
  wire [7:0] R0_data_0_58 = mem_0_58_R0_data;
  wire [7:0] R0_data_0_59 = mem_0_59_R0_data;
  wire [7:0] R0_data_0_60 = mem_0_60_R0_data;
  wire [7:0] R0_data_0_61 = mem_0_61_R0_data;
  wire [7:0] R0_data_0_62 = mem_0_62_R0_data;
  wire [7:0] R0_data_0_63 = mem_0_63_R0_data;
  wire [15:0] _GEN_0 = {R0_data_0_1,R0_data_0_0};
  wire [23:0] _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [31:0] _GEN_2 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [39:0] _GEN_3 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [47:0] _GEN_4 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [55:0] _GEN_5 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [63:0] _GEN_6 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}
    ;
  wire [71:0] _GEN_7 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,
    R0_data_0_0};
  wire [79:0] _GEN_8 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,
    R0_data_0_1,R0_data_0_0};
  wire [87:0] _GEN_9 = {R0_data_0_10,_GEN_8};
  wire [95:0] _GEN_10 = {R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [103:0] _GEN_11 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [111:0] _GEN_12 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [119:0] _GEN_13 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [127:0] _GEN_14 = {R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [135:0] _GEN_15 = {R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,
    _GEN_8};
  wire [143:0] _GEN_16 = {R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,
    R0_data_0_10,_GEN_8};
  wire [151:0] _GEN_17 = {R0_data_0_18,R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,
    R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [159:0] _GEN_18 = {R0_data_0_19,_GEN_17};
  wire [167:0] _GEN_19 = {R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [175:0] _GEN_20 = {R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [183:0] _GEN_21 = {R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [191:0] _GEN_22 = {R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [199:0] _GEN_23 = {R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [207:0] _GEN_24 = {R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,
    _GEN_17};
  wire [215:0] _GEN_25 = {R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,
    R0_data_0_19,_GEN_17};
  wire [223:0] _GEN_26 = {R0_data_0_27,R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,
    R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [231:0] _GEN_27 = {R0_data_0_28,_GEN_26};
  wire [239:0] _GEN_28 = {R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [247:0] _GEN_29 = {R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [255:0] _GEN_30 = {R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [263:0] _GEN_31 = {R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [271:0] _GEN_32 = {R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [279:0] _GEN_33 = {R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,
    _GEN_26};
  wire [287:0] _GEN_34 = {R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,
    R0_data_0_28,_GEN_26};
  wire [295:0] _GEN_35 = {R0_data_0_36,R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,
    R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [303:0] _GEN_36 = {R0_data_0_37,_GEN_35};
  wire [311:0] _GEN_37 = {R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [319:0] _GEN_38 = {R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [327:0] _GEN_39 = {R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [335:0] _GEN_40 = {R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [343:0] _GEN_41 = {R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [351:0] _GEN_42 = {R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,
    _GEN_35};
  wire [359:0] _GEN_43 = {R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,
    R0_data_0_37,_GEN_35};
  wire [367:0] _GEN_44 = {R0_data_0_45,R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,
    R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [375:0] _GEN_45 = {R0_data_0_46,_GEN_44};
  wire [383:0] _GEN_46 = {R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [391:0] _GEN_47 = {R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [399:0] _GEN_48 = {R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [407:0] _GEN_49 = {R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [415:0] _GEN_50 = {R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [423:0] _GEN_51 = {R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,
    _GEN_44};
  wire [431:0] _GEN_52 = {R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,
    R0_data_0_46,_GEN_44};
  wire [439:0] _GEN_53 = {R0_data_0_54,R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,
    R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [447:0] _GEN_54 = {R0_data_0_55,_GEN_53};
  wire [455:0] _GEN_55 = {R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [463:0] _GEN_56 = {R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [471:0] _GEN_57 = {R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [479:0] _GEN_58 = {R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [487:0] _GEN_59 = {R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [495:0] _GEN_60 = {R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,
    _GEN_53};
  wire [503:0] _GEN_61 = {R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,
    R0_data_0_55,_GEN_53};
  wire [511:0] R0_data_0 = {R0_data_0_63,R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,
    R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [15:0] _GEN_62 = {R0_data_0_1,R0_data_0_0};
  wire [23:0] _GEN_63 = {R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [31:0] _GEN_64 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [39:0] _GEN_65 = {R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [47:0] _GEN_66 = {R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [55:0] _GEN_67 = {R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [63:0] _GEN_68 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0
    };
  wire [71:0] _GEN_69 = {R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1
    ,R0_data_0_0};
  wire [79:0] _GEN_70 = {R0_data_0_9,R0_data_0_8,R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2
    ,R0_data_0_1,R0_data_0_0};
  wire [87:0] _GEN_71 = {R0_data_0_10,_GEN_8};
  wire [95:0] _GEN_72 = {R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [103:0] _GEN_73 = {R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [111:0] _GEN_74 = {R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [119:0] _GEN_75 = {R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [127:0] _GEN_76 = {R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [135:0] _GEN_77 = {R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,R0_data_0_10,
    _GEN_8};
  wire [143:0] _GEN_78 = {R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,R0_data_0_11,
    R0_data_0_10,_GEN_8};
  wire [151:0] _GEN_79 = {R0_data_0_18,R0_data_0_17,R0_data_0_16,R0_data_0_15,R0_data_0_14,R0_data_0_13,R0_data_0_12,
    R0_data_0_11,R0_data_0_10,_GEN_8};
  wire [159:0] _GEN_80 = {R0_data_0_19,_GEN_17};
  wire [167:0] _GEN_81 = {R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [175:0] _GEN_82 = {R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [183:0] _GEN_83 = {R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [191:0] _GEN_84 = {R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [199:0] _GEN_85 = {R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [207:0] _GEN_86 = {R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,R0_data_0_19,
    _GEN_17};
  wire [215:0] _GEN_87 = {R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,R0_data_0_20,
    R0_data_0_19,_GEN_17};
  wire [223:0] _GEN_88 = {R0_data_0_27,R0_data_0_26,R0_data_0_25,R0_data_0_24,R0_data_0_23,R0_data_0_22,R0_data_0_21,
    R0_data_0_20,R0_data_0_19,_GEN_17};
  wire [231:0] _GEN_89 = {R0_data_0_28,_GEN_26};
  wire [239:0] _GEN_90 = {R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [247:0] _GEN_91 = {R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [255:0] _GEN_92 = {R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [263:0] _GEN_93 = {R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [271:0] _GEN_94 = {R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [279:0] _GEN_95 = {R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,R0_data_0_28,
    _GEN_26};
  wire [287:0] _GEN_96 = {R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,R0_data_0_29,
    R0_data_0_28,_GEN_26};
  wire [295:0] _GEN_97 = {R0_data_0_36,R0_data_0_35,R0_data_0_34,R0_data_0_33,R0_data_0_32,R0_data_0_31,R0_data_0_30,
    R0_data_0_29,R0_data_0_28,_GEN_26};
  wire [303:0] _GEN_98 = {R0_data_0_37,_GEN_35};
  wire [311:0] _GEN_99 = {R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [319:0] _GEN_100 = {R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [327:0] _GEN_101 = {R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [335:0] _GEN_102 = {R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [343:0] _GEN_103 = {R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [351:0] _GEN_104 = {R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,R0_data_0_37,
    _GEN_35};
  wire [359:0] _GEN_105 = {R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,R0_data_0_38,
    R0_data_0_37,_GEN_35};
  wire [367:0] _GEN_106 = {R0_data_0_45,R0_data_0_44,R0_data_0_43,R0_data_0_42,R0_data_0_41,R0_data_0_40,R0_data_0_39,
    R0_data_0_38,R0_data_0_37,_GEN_35};
  wire [375:0] _GEN_107 = {R0_data_0_46,_GEN_44};
  wire [383:0] _GEN_108 = {R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [391:0] _GEN_109 = {R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [399:0] _GEN_110 = {R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [407:0] _GEN_111 = {R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [415:0] _GEN_112 = {R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [423:0] _GEN_113 = {R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,R0_data_0_46,
    _GEN_44};
  wire [431:0] _GEN_114 = {R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,R0_data_0_47,
    R0_data_0_46,_GEN_44};
  wire [439:0] _GEN_115 = {R0_data_0_54,R0_data_0_53,R0_data_0_52,R0_data_0_51,R0_data_0_50,R0_data_0_49,R0_data_0_48,
    R0_data_0_47,R0_data_0_46,_GEN_44};
  wire [447:0] _GEN_116 = {R0_data_0_55,_GEN_53};
  wire [455:0] _GEN_117 = {R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [463:0] _GEN_118 = {R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [471:0] _GEN_119 = {R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [479:0] _GEN_120 = {R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [487:0] _GEN_121 = {R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,_GEN_53};
  wire [495:0] _GEN_122 = {R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,R0_data_0_55,
    _GEN_53};
  wire [503:0] _GEN_123 = {R0_data_0_62,R0_data_0_61,R0_data_0_60,R0_data_0_59,R0_data_0_58,R0_data_0_57,R0_data_0_56,
    R0_data_0_55,_GEN_53};
  split_mem_0_ext mem_0_0 (
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en),
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask)
  );
  split_mem_0_ext mem_0_1 (
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en),
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask)
  );
  split_mem_0_ext mem_0_2 (
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en),
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask)
  );
  split_mem_0_ext mem_0_3 (
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en),
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask)
  );
  split_mem_0_ext mem_0_4 (
    .R0_addr(mem_0_4_R0_addr),
    .R0_clk(mem_0_4_R0_clk),
    .R0_data(mem_0_4_R0_data),
    .R0_en(mem_0_4_R0_en),
    .W0_addr(mem_0_4_W0_addr),
    .W0_clk(mem_0_4_W0_clk),
    .W0_data(mem_0_4_W0_data),
    .W0_en(mem_0_4_W0_en),
    .W0_mask(mem_0_4_W0_mask)
  );
  split_mem_0_ext mem_0_5 (
    .R0_addr(mem_0_5_R0_addr),
    .R0_clk(mem_0_5_R0_clk),
    .R0_data(mem_0_5_R0_data),
    .R0_en(mem_0_5_R0_en),
    .W0_addr(mem_0_5_W0_addr),
    .W0_clk(mem_0_5_W0_clk),
    .W0_data(mem_0_5_W0_data),
    .W0_en(mem_0_5_W0_en),
    .W0_mask(mem_0_5_W0_mask)
  );
  split_mem_0_ext mem_0_6 (
    .R0_addr(mem_0_6_R0_addr),
    .R0_clk(mem_0_6_R0_clk),
    .R0_data(mem_0_6_R0_data),
    .R0_en(mem_0_6_R0_en),
    .W0_addr(mem_0_6_W0_addr),
    .W0_clk(mem_0_6_W0_clk),
    .W0_data(mem_0_6_W0_data),
    .W0_en(mem_0_6_W0_en),
    .W0_mask(mem_0_6_W0_mask)
  );
  split_mem_0_ext mem_0_7 (
    .R0_addr(mem_0_7_R0_addr),
    .R0_clk(mem_0_7_R0_clk),
    .R0_data(mem_0_7_R0_data),
    .R0_en(mem_0_7_R0_en),
    .W0_addr(mem_0_7_W0_addr),
    .W0_clk(mem_0_7_W0_clk),
    .W0_data(mem_0_7_W0_data),
    .W0_en(mem_0_7_W0_en),
    .W0_mask(mem_0_7_W0_mask)
  );
  split_mem_0_ext mem_0_8 (
    .R0_addr(mem_0_8_R0_addr),
    .R0_clk(mem_0_8_R0_clk),
    .R0_data(mem_0_8_R0_data),
    .R0_en(mem_0_8_R0_en),
    .W0_addr(mem_0_8_W0_addr),
    .W0_clk(mem_0_8_W0_clk),
    .W0_data(mem_0_8_W0_data),
    .W0_en(mem_0_8_W0_en),
    .W0_mask(mem_0_8_W0_mask)
  );
  split_mem_0_ext mem_0_9 (
    .R0_addr(mem_0_9_R0_addr),
    .R0_clk(mem_0_9_R0_clk),
    .R0_data(mem_0_9_R0_data),
    .R0_en(mem_0_9_R0_en),
    .W0_addr(mem_0_9_W0_addr),
    .W0_clk(mem_0_9_W0_clk),
    .W0_data(mem_0_9_W0_data),
    .W0_en(mem_0_9_W0_en),
    .W0_mask(mem_0_9_W0_mask)
  );
  split_mem_0_ext mem_0_10 (
    .R0_addr(mem_0_10_R0_addr),
    .R0_clk(mem_0_10_R0_clk),
    .R0_data(mem_0_10_R0_data),
    .R0_en(mem_0_10_R0_en),
    .W0_addr(mem_0_10_W0_addr),
    .W0_clk(mem_0_10_W0_clk),
    .W0_data(mem_0_10_W0_data),
    .W0_en(mem_0_10_W0_en),
    .W0_mask(mem_0_10_W0_mask)
  );
  split_mem_0_ext mem_0_11 (
    .R0_addr(mem_0_11_R0_addr),
    .R0_clk(mem_0_11_R0_clk),
    .R0_data(mem_0_11_R0_data),
    .R0_en(mem_0_11_R0_en),
    .W0_addr(mem_0_11_W0_addr),
    .W0_clk(mem_0_11_W0_clk),
    .W0_data(mem_0_11_W0_data),
    .W0_en(mem_0_11_W0_en),
    .W0_mask(mem_0_11_W0_mask)
  );
  split_mem_0_ext mem_0_12 (
    .R0_addr(mem_0_12_R0_addr),
    .R0_clk(mem_0_12_R0_clk),
    .R0_data(mem_0_12_R0_data),
    .R0_en(mem_0_12_R0_en),
    .W0_addr(mem_0_12_W0_addr),
    .W0_clk(mem_0_12_W0_clk),
    .W0_data(mem_0_12_W0_data),
    .W0_en(mem_0_12_W0_en),
    .W0_mask(mem_0_12_W0_mask)
  );
  split_mem_0_ext mem_0_13 (
    .R0_addr(mem_0_13_R0_addr),
    .R0_clk(mem_0_13_R0_clk),
    .R0_data(mem_0_13_R0_data),
    .R0_en(mem_0_13_R0_en),
    .W0_addr(mem_0_13_W0_addr),
    .W0_clk(mem_0_13_W0_clk),
    .W0_data(mem_0_13_W0_data),
    .W0_en(mem_0_13_W0_en),
    .W0_mask(mem_0_13_W0_mask)
  );
  split_mem_0_ext mem_0_14 (
    .R0_addr(mem_0_14_R0_addr),
    .R0_clk(mem_0_14_R0_clk),
    .R0_data(mem_0_14_R0_data),
    .R0_en(mem_0_14_R0_en),
    .W0_addr(mem_0_14_W0_addr),
    .W0_clk(mem_0_14_W0_clk),
    .W0_data(mem_0_14_W0_data),
    .W0_en(mem_0_14_W0_en),
    .W0_mask(mem_0_14_W0_mask)
  );
  split_mem_0_ext mem_0_15 (
    .R0_addr(mem_0_15_R0_addr),
    .R0_clk(mem_0_15_R0_clk),
    .R0_data(mem_0_15_R0_data),
    .R0_en(mem_0_15_R0_en),
    .W0_addr(mem_0_15_W0_addr),
    .W0_clk(mem_0_15_W0_clk),
    .W0_data(mem_0_15_W0_data),
    .W0_en(mem_0_15_W0_en),
    .W0_mask(mem_0_15_W0_mask)
  );
  split_mem_0_ext mem_0_16 (
    .R0_addr(mem_0_16_R0_addr),
    .R0_clk(mem_0_16_R0_clk),
    .R0_data(mem_0_16_R0_data),
    .R0_en(mem_0_16_R0_en),
    .W0_addr(mem_0_16_W0_addr),
    .W0_clk(mem_0_16_W0_clk),
    .W0_data(mem_0_16_W0_data),
    .W0_en(mem_0_16_W0_en),
    .W0_mask(mem_0_16_W0_mask)
  );
  split_mem_0_ext mem_0_17 (
    .R0_addr(mem_0_17_R0_addr),
    .R0_clk(mem_0_17_R0_clk),
    .R0_data(mem_0_17_R0_data),
    .R0_en(mem_0_17_R0_en),
    .W0_addr(mem_0_17_W0_addr),
    .W0_clk(mem_0_17_W0_clk),
    .W0_data(mem_0_17_W0_data),
    .W0_en(mem_0_17_W0_en),
    .W0_mask(mem_0_17_W0_mask)
  );
  split_mem_0_ext mem_0_18 (
    .R0_addr(mem_0_18_R0_addr),
    .R0_clk(mem_0_18_R0_clk),
    .R0_data(mem_0_18_R0_data),
    .R0_en(mem_0_18_R0_en),
    .W0_addr(mem_0_18_W0_addr),
    .W0_clk(mem_0_18_W0_clk),
    .W0_data(mem_0_18_W0_data),
    .W0_en(mem_0_18_W0_en),
    .W0_mask(mem_0_18_W0_mask)
  );
  split_mem_0_ext mem_0_19 (
    .R0_addr(mem_0_19_R0_addr),
    .R0_clk(mem_0_19_R0_clk),
    .R0_data(mem_0_19_R0_data),
    .R0_en(mem_0_19_R0_en),
    .W0_addr(mem_0_19_W0_addr),
    .W0_clk(mem_0_19_W0_clk),
    .W0_data(mem_0_19_W0_data),
    .W0_en(mem_0_19_W0_en),
    .W0_mask(mem_0_19_W0_mask)
  );
  split_mem_0_ext mem_0_20 (
    .R0_addr(mem_0_20_R0_addr),
    .R0_clk(mem_0_20_R0_clk),
    .R0_data(mem_0_20_R0_data),
    .R0_en(mem_0_20_R0_en),
    .W0_addr(mem_0_20_W0_addr),
    .W0_clk(mem_0_20_W0_clk),
    .W0_data(mem_0_20_W0_data),
    .W0_en(mem_0_20_W0_en),
    .W0_mask(mem_0_20_W0_mask)
  );
  split_mem_0_ext mem_0_21 (
    .R0_addr(mem_0_21_R0_addr),
    .R0_clk(mem_0_21_R0_clk),
    .R0_data(mem_0_21_R0_data),
    .R0_en(mem_0_21_R0_en),
    .W0_addr(mem_0_21_W0_addr),
    .W0_clk(mem_0_21_W0_clk),
    .W0_data(mem_0_21_W0_data),
    .W0_en(mem_0_21_W0_en),
    .W0_mask(mem_0_21_W0_mask)
  );
  split_mem_0_ext mem_0_22 (
    .R0_addr(mem_0_22_R0_addr),
    .R0_clk(mem_0_22_R0_clk),
    .R0_data(mem_0_22_R0_data),
    .R0_en(mem_0_22_R0_en),
    .W0_addr(mem_0_22_W0_addr),
    .W0_clk(mem_0_22_W0_clk),
    .W0_data(mem_0_22_W0_data),
    .W0_en(mem_0_22_W0_en),
    .W0_mask(mem_0_22_W0_mask)
  );
  split_mem_0_ext mem_0_23 (
    .R0_addr(mem_0_23_R0_addr),
    .R0_clk(mem_0_23_R0_clk),
    .R0_data(mem_0_23_R0_data),
    .R0_en(mem_0_23_R0_en),
    .W0_addr(mem_0_23_W0_addr),
    .W0_clk(mem_0_23_W0_clk),
    .W0_data(mem_0_23_W0_data),
    .W0_en(mem_0_23_W0_en),
    .W0_mask(mem_0_23_W0_mask)
  );
  split_mem_0_ext mem_0_24 (
    .R0_addr(mem_0_24_R0_addr),
    .R0_clk(mem_0_24_R0_clk),
    .R0_data(mem_0_24_R0_data),
    .R0_en(mem_0_24_R0_en),
    .W0_addr(mem_0_24_W0_addr),
    .W0_clk(mem_0_24_W0_clk),
    .W0_data(mem_0_24_W0_data),
    .W0_en(mem_0_24_W0_en),
    .W0_mask(mem_0_24_W0_mask)
  );
  split_mem_0_ext mem_0_25 (
    .R0_addr(mem_0_25_R0_addr),
    .R0_clk(mem_0_25_R0_clk),
    .R0_data(mem_0_25_R0_data),
    .R0_en(mem_0_25_R0_en),
    .W0_addr(mem_0_25_W0_addr),
    .W0_clk(mem_0_25_W0_clk),
    .W0_data(mem_0_25_W0_data),
    .W0_en(mem_0_25_W0_en),
    .W0_mask(mem_0_25_W0_mask)
  );
  split_mem_0_ext mem_0_26 (
    .R0_addr(mem_0_26_R0_addr),
    .R0_clk(mem_0_26_R0_clk),
    .R0_data(mem_0_26_R0_data),
    .R0_en(mem_0_26_R0_en),
    .W0_addr(mem_0_26_W0_addr),
    .W0_clk(mem_0_26_W0_clk),
    .W0_data(mem_0_26_W0_data),
    .W0_en(mem_0_26_W0_en),
    .W0_mask(mem_0_26_W0_mask)
  );
  split_mem_0_ext mem_0_27 (
    .R0_addr(mem_0_27_R0_addr),
    .R0_clk(mem_0_27_R0_clk),
    .R0_data(mem_0_27_R0_data),
    .R0_en(mem_0_27_R0_en),
    .W0_addr(mem_0_27_W0_addr),
    .W0_clk(mem_0_27_W0_clk),
    .W0_data(mem_0_27_W0_data),
    .W0_en(mem_0_27_W0_en),
    .W0_mask(mem_0_27_W0_mask)
  );
  split_mem_0_ext mem_0_28 (
    .R0_addr(mem_0_28_R0_addr),
    .R0_clk(mem_0_28_R0_clk),
    .R0_data(mem_0_28_R0_data),
    .R0_en(mem_0_28_R0_en),
    .W0_addr(mem_0_28_W0_addr),
    .W0_clk(mem_0_28_W0_clk),
    .W0_data(mem_0_28_W0_data),
    .W0_en(mem_0_28_W0_en),
    .W0_mask(mem_0_28_W0_mask)
  );
  split_mem_0_ext mem_0_29 (
    .R0_addr(mem_0_29_R0_addr),
    .R0_clk(mem_0_29_R0_clk),
    .R0_data(mem_0_29_R0_data),
    .R0_en(mem_0_29_R0_en),
    .W0_addr(mem_0_29_W0_addr),
    .W0_clk(mem_0_29_W0_clk),
    .W0_data(mem_0_29_W0_data),
    .W0_en(mem_0_29_W0_en),
    .W0_mask(mem_0_29_W0_mask)
  );
  split_mem_0_ext mem_0_30 (
    .R0_addr(mem_0_30_R0_addr),
    .R0_clk(mem_0_30_R0_clk),
    .R0_data(mem_0_30_R0_data),
    .R0_en(mem_0_30_R0_en),
    .W0_addr(mem_0_30_W0_addr),
    .W0_clk(mem_0_30_W0_clk),
    .W0_data(mem_0_30_W0_data),
    .W0_en(mem_0_30_W0_en),
    .W0_mask(mem_0_30_W0_mask)
  );
  split_mem_0_ext mem_0_31 (
    .R0_addr(mem_0_31_R0_addr),
    .R0_clk(mem_0_31_R0_clk),
    .R0_data(mem_0_31_R0_data),
    .R0_en(mem_0_31_R0_en),
    .W0_addr(mem_0_31_W0_addr),
    .W0_clk(mem_0_31_W0_clk),
    .W0_data(mem_0_31_W0_data),
    .W0_en(mem_0_31_W0_en),
    .W0_mask(mem_0_31_W0_mask)
  );
  split_mem_0_ext mem_0_32 (
    .R0_addr(mem_0_32_R0_addr),
    .R0_clk(mem_0_32_R0_clk),
    .R0_data(mem_0_32_R0_data),
    .R0_en(mem_0_32_R0_en),
    .W0_addr(mem_0_32_W0_addr),
    .W0_clk(mem_0_32_W0_clk),
    .W0_data(mem_0_32_W0_data),
    .W0_en(mem_0_32_W0_en),
    .W0_mask(mem_0_32_W0_mask)
  );
  split_mem_0_ext mem_0_33 (
    .R0_addr(mem_0_33_R0_addr),
    .R0_clk(mem_0_33_R0_clk),
    .R0_data(mem_0_33_R0_data),
    .R0_en(mem_0_33_R0_en),
    .W0_addr(mem_0_33_W0_addr),
    .W0_clk(mem_0_33_W0_clk),
    .W0_data(mem_0_33_W0_data),
    .W0_en(mem_0_33_W0_en),
    .W0_mask(mem_0_33_W0_mask)
  );
  split_mem_0_ext mem_0_34 (
    .R0_addr(mem_0_34_R0_addr),
    .R0_clk(mem_0_34_R0_clk),
    .R0_data(mem_0_34_R0_data),
    .R0_en(mem_0_34_R0_en),
    .W0_addr(mem_0_34_W0_addr),
    .W0_clk(mem_0_34_W0_clk),
    .W0_data(mem_0_34_W0_data),
    .W0_en(mem_0_34_W0_en),
    .W0_mask(mem_0_34_W0_mask)
  );
  split_mem_0_ext mem_0_35 (
    .R0_addr(mem_0_35_R0_addr),
    .R0_clk(mem_0_35_R0_clk),
    .R0_data(mem_0_35_R0_data),
    .R0_en(mem_0_35_R0_en),
    .W0_addr(mem_0_35_W0_addr),
    .W0_clk(mem_0_35_W0_clk),
    .W0_data(mem_0_35_W0_data),
    .W0_en(mem_0_35_W0_en),
    .W0_mask(mem_0_35_W0_mask)
  );
  split_mem_0_ext mem_0_36 (
    .R0_addr(mem_0_36_R0_addr),
    .R0_clk(mem_0_36_R0_clk),
    .R0_data(mem_0_36_R0_data),
    .R0_en(mem_0_36_R0_en),
    .W0_addr(mem_0_36_W0_addr),
    .W0_clk(mem_0_36_W0_clk),
    .W0_data(mem_0_36_W0_data),
    .W0_en(mem_0_36_W0_en),
    .W0_mask(mem_0_36_W0_mask)
  );
  split_mem_0_ext mem_0_37 (
    .R0_addr(mem_0_37_R0_addr),
    .R0_clk(mem_0_37_R0_clk),
    .R0_data(mem_0_37_R0_data),
    .R0_en(mem_0_37_R0_en),
    .W0_addr(mem_0_37_W0_addr),
    .W0_clk(mem_0_37_W0_clk),
    .W0_data(mem_0_37_W0_data),
    .W0_en(mem_0_37_W0_en),
    .W0_mask(mem_0_37_W0_mask)
  );
  split_mem_0_ext mem_0_38 (
    .R0_addr(mem_0_38_R0_addr),
    .R0_clk(mem_0_38_R0_clk),
    .R0_data(mem_0_38_R0_data),
    .R0_en(mem_0_38_R0_en),
    .W0_addr(mem_0_38_W0_addr),
    .W0_clk(mem_0_38_W0_clk),
    .W0_data(mem_0_38_W0_data),
    .W0_en(mem_0_38_W0_en),
    .W0_mask(mem_0_38_W0_mask)
  );
  split_mem_0_ext mem_0_39 (
    .R0_addr(mem_0_39_R0_addr),
    .R0_clk(mem_0_39_R0_clk),
    .R0_data(mem_0_39_R0_data),
    .R0_en(mem_0_39_R0_en),
    .W0_addr(mem_0_39_W0_addr),
    .W0_clk(mem_0_39_W0_clk),
    .W0_data(mem_0_39_W0_data),
    .W0_en(mem_0_39_W0_en),
    .W0_mask(mem_0_39_W0_mask)
  );
  split_mem_0_ext mem_0_40 (
    .R0_addr(mem_0_40_R0_addr),
    .R0_clk(mem_0_40_R0_clk),
    .R0_data(mem_0_40_R0_data),
    .R0_en(mem_0_40_R0_en),
    .W0_addr(mem_0_40_W0_addr),
    .W0_clk(mem_0_40_W0_clk),
    .W0_data(mem_0_40_W0_data),
    .W0_en(mem_0_40_W0_en),
    .W0_mask(mem_0_40_W0_mask)
  );
  split_mem_0_ext mem_0_41 (
    .R0_addr(mem_0_41_R0_addr),
    .R0_clk(mem_0_41_R0_clk),
    .R0_data(mem_0_41_R0_data),
    .R0_en(mem_0_41_R0_en),
    .W0_addr(mem_0_41_W0_addr),
    .W0_clk(mem_0_41_W0_clk),
    .W0_data(mem_0_41_W0_data),
    .W0_en(mem_0_41_W0_en),
    .W0_mask(mem_0_41_W0_mask)
  );
  split_mem_0_ext mem_0_42 (
    .R0_addr(mem_0_42_R0_addr),
    .R0_clk(mem_0_42_R0_clk),
    .R0_data(mem_0_42_R0_data),
    .R0_en(mem_0_42_R0_en),
    .W0_addr(mem_0_42_W0_addr),
    .W0_clk(mem_0_42_W0_clk),
    .W0_data(mem_0_42_W0_data),
    .W0_en(mem_0_42_W0_en),
    .W0_mask(mem_0_42_W0_mask)
  );
  split_mem_0_ext mem_0_43 (
    .R0_addr(mem_0_43_R0_addr),
    .R0_clk(mem_0_43_R0_clk),
    .R0_data(mem_0_43_R0_data),
    .R0_en(mem_0_43_R0_en),
    .W0_addr(mem_0_43_W0_addr),
    .W0_clk(mem_0_43_W0_clk),
    .W0_data(mem_0_43_W0_data),
    .W0_en(mem_0_43_W0_en),
    .W0_mask(mem_0_43_W0_mask)
  );
  split_mem_0_ext mem_0_44 (
    .R0_addr(mem_0_44_R0_addr),
    .R0_clk(mem_0_44_R0_clk),
    .R0_data(mem_0_44_R0_data),
    .R0_en(mem_0_44_R0_en),
    .W0_addr(mem_0_44_W0_addr),
    .W0_clk(mem_0_44_W0_clk),
    .W0_data(mem_0_44_W0_data),
    .W0_en(mem_0_44_W0_en),
    .W0_mask(mem_0_44_W0_mask)
  );
  split_mem_0_ext mem_0_45 (
    .R0_addr(mem_0_45_R0_addr),
    .R0_clk(mem_0_45_R0_clk),
    .R0_data(mem_0_45_R0_data),
    .R0_en(mem_0_45_R0_en),
    .W0_addr(mem_0_45_W0_addr),
    .W0_clk(mem_0_45_W0_clk),
    .W0_data(mem_0_45_W0_data),
    .W0_en(mem_0_45_W0_en),
    .W0_mask(mem_0_45_W0_mask)
  );
  split_mem_0_ext mem_0_46 (
    .R0_addr(mem_0_46_R0_addr),
    .R0_clk(mem_0_46_R0_clk),
    .R0_data(mem_0_46_R0_data),
    .R0_en(mem_0_46_R0_en),
    .W0_addr(mem_0_46_W0_addr),
    .W0_clk(mem_0_46_W0_clk),
    .W0_data(mem_0_46_W0_data),
    .W0_en(mem_0_46_W0_en),
    .W0_mask(mem_0_46_W0_mask)
  );
  split_mem_0_ext mem_0_47 (
    .R0_addr(mem_0_47_R0_addr),
    .R0_clk(mem_0_47_R0_clk),
    .R0_data(mem_0_47_R0_data),
    .R0_en(mem_0_47_R0_en),
    .W0_addr(mem_0_47_W0_addr),
    .W0_clk(mem_0_47_W0_clk),
    .W0_data(mem_0_47_W0_data),
    .W0_en(mem_0_47_W0_en),
    .W0_mask(mem_0_47_W0_mask)
  );
  split_mem_0_ext mem_0_48 (
    .R0_addr(mem_0_48_R0_addr),
    .R0_clk(mem_0_48_R0_clk),
    .R0_data(mem_0_48_R0_data),
    .R0_en(mem_0_48_R0_en),
    .W0_addr(mem_0_48_W0_addr),
    .W0_clk(mem_0_48_W0_clk),
    .W0_data(mem_0_48_W0_data),
    .W0_en(mem_0_48_W0_en),
    .W0_mask(mem_0_48_W0_mask)
  );
  split_mem_0_ext mem_0_49 (
    .R0_addr(mem_0_49_R0_addr),
    .R0_clk(mem_0_49_R0_clk),
    .R0_data(mem_0_49_R0_data),
    .R0_en(mem_0_49_R0_en),
    .W0_addr(mem_0_49_W0_addr),
    .W0_clk(mem_0_49_W0_clk),
    .W0_data(mem_0_49_W0_data),
    .W0_en(mem_0_49_W0_en),
    .W0_mask(mem_0_49_W0_mask)
  );
  split_mem_0_ext mem_0_50 (
    .R0_addr(mem_0_50_R0_addr),
    .R0_clk(mem_0_50_R0_clk),
    .R0_data(mem_0_50_R0_data),
    .R0_en(mem_0_50_R0_en),
    .W0_addr(mem_0_50_W0_addr),
    .W0_clk(mem_0_50_W0_clk),
    .W0_data(mem_0_50_W0_data),
    .W0_en(mem_0_50_W0_en),
    .W0_mask(mem_0_50_W0_mask)
  );
  split_mem_0_ext mem_0_51 (
    .R0_addr(mem_0_51_R0_addr),
    .R0_clk(mem_0_51_R0_clk),
    .R0_data(mem_0_51_R0_data),
    .R0_en(mem_0_51_R0_en),
    .W0_addr(mem_0_51_W0_addr),
    .W0_clk(mem_0_51_W0_clk),
    .W0_data(mem_0_51_W0_data),
    .W0_en(mem_0_51_W0_en),
    .W0_mask(mem_0_51_W0_mask)
  );
  split_mem_0_ext mem_0_52 (
    .R0_addr(mem_0_52_R0_addr),
    .R0_clk(mem_0_52_R0_clk),
    .R0_data(mem_0_52_R0_data),
    .R0_en(mem_0_52_R0_en),
    .W0_addr(mem_0_52_W0_addr),
    .W0_clk(mem_0_52_W0_clk),
    .W0_data(mem_0_52_W0_data),
    .W0_en(mem_0_52_W0_en),
    .W0_mask(mem_0_52_W0_mask)
  );
  split_mem_0_ext mem_0_53 (
    .R0_addr(mem_0_53_R0_addr),
    .R0_clk(mem_0_53_R0_clk),
    .R0_data(mem_0_53_R0_data),
    .R0_en(mem_0_53_R0_en),
    .W0_addr(mem_0_53_W0_addr),
    .W0_clk(mem_0_53_W0_clk),
    .W0_data(mem_0_53_W0_data),
    .W0_en(mem_0_53_W0_en),
    .W0_mask(mem_0_53_W0_mask)
  );
  split_mem_0_ext mem_0_54 (
    .R0_addr(mem_0_54_R0_addr),
    .R0_clk(mem_0_54_R0_clk),
    .R0_data(mem_0_54_R0_data),
    .R0_en(mem_0_54_R0_en),
    .W0_addr(mem_0_54_W0_addr),
    .W0_clk(mem_0_54_W0_clk),
    .W0_data(mem_0_54_W0_data),
    .W0_en(mem_0_54_W0_en),
    .W0_mask(mem_0_54_W0_mask)
  );
  split_mem_0_ext mem_0_55 (
    .R0_addr(mem_0_55_R0_addr),
    .R0_clk(mem_0_55_R0_clk),
    .R0_data(mem_0_55_R0_data),
    .R0_en(mem_0_55_R0_en),
    .W0_addr(mem_0_55_W0_addr),
    .W0_clk(mem_0_55_W0_clk),
    .W0_data(mem_0_55_W0_data),
    .W0_en(mem_0_55_W0_en),
    .W0_mask(mem_0_55_W0_mask)
  );
  split_mem_0_ext mem_0_56 (
    .R0_addr(mem_0_56_R0_addr),
    .R0_clk(mem_0_56_R0_clk),
    .R0_data(mem_0_56_R0_data),
    .R0_en(mem_0_56_R0_en),
    .W0_addr(mem_0_56_W0_addr),
    .W0_clk(mem_0_56_W0_clk),
    .W0_data(mem_0_56_W0_data),
    .W0_en(mem_0_56_W0_en),
    .W0_mask(mem_0_56_W0_mask)
  );
  split_mem_0_ext mem_0_57 (
    .R0_addr(mem_0_57_R0_addr),
    .R0_clk(mem_0_57_R0_clk),
    .R0_data(mem_0_57_R0_data),
    .R0_en(mem_0_57_R0_en),
    .W0_addr(mem_0_57_W0_addr),
    .W0_clk(mem_0_57_W0_clk),
    .W0_data(mem_0_57_W0_data),
    .W0_en(mem_0_57_W0_en),
    .W0_mask(mem_0_57_W0_mask)
  );
  split_mem_0_ext mem_0_58 (
    .R0_addr(mem_0_58_R0_addr),
    .R0_clk(mem_0_58_R0_clk),
    .R0_data(mem_0_58_R0_data),
    .R0_en(mem_0_58_R0_en),
    .W0_addr(mem_0_58_W0_addr),
    .W0_clk(mem_0_58_W0_clk),
    .W0_data(mem_0_58_W0_data),
    .W0_en(mem_0_58_W0_en),
    .W0_mask(mem_0_58_W0_mask)
  );
  split_mem_0_ext mem_0_59 (
    .R0_addr(mem_0_59_R0_addr),
    .R0_clk(mem_0_59_R0_clk),
    .R0_data(mem_0_59_R0_data),
    .R0_en(mem_0_59_R0_en),
    .W0_addr(mem_0_59_W0_addr),
    .W0_clk(mem_0_59_W0_clk),
    .W0_data(mem_0_59_W0_data),
    .W0_en(mem_0_59_W0_en),
    .W0_mask(mem_0_59_W0_mask)
  );
  split_mem_0_ext mem_0_60 (
    .R0_addr(mem_0_60_R0_addr),
    .R0_clk(mem_0_60_R0_clk),
    .R0_data(mem_0_60_R0_data),
    .R0_en(mem_0_60_R0_en),
    .W0_addr(mem_0_60_W0_addr),
    .W0_clk(mem_0_60_W0_clk),
    .W0_data(mem_0_60_W0_data),
    .W0_en(mem_0_60_W0_en),
    .W0_mask(mem_0_60_W0_mask)
  );
  split_mem_0_ext mem_0_61 (
    .R0_addr(mem_0_61_R0_addr),
    .R0_clk(mem_0_61_R0_clk),
    .R0_data(mem_0_61_R0_data),
    .R0_en(mem_0_61_R0_en),
    .W0_addr(mem_0_61_W0_addr),
    .W0_clk(mem_0_61_W0_clk),
    .W0_data(mem_0_61_W0_data),
    .W0_en(mem_0_61_W0_en),
    .W0_mask(mem_0_61_W0_mask)
  );
  split_mem_0_ext mem_0_62 (
    .R0_addr(mem_0_62_R0_addr),
    .R0_clk(mem_0_62_R0_clk),
    .R0_data(mem_0_62_R0_data),
    .R0_en(mem_0_62_R0_en),
    .W0_addr(mem_0_62_W0_addr),
    .W0_clk(mem_0_62_W0_clk),
    .W0_data(mem_0_62_W0_data),
    .W0_en(mem_0_62_W0_en),
    .W0_mask(mem_0_62_W0_mask)
  );
  split_mem_0_ext mem_0_63 (
    .R0_addr(mem_0_63_R0_addr),
    .R0_clk(mem_0_63_R0_clk),
    .R0_data(mem_0_63_R0_data),
    .R0_en(mem_0_63_R0_en),
    .W0_addr(mem_0_63_W0_addr),
    .W0_clk(mem_0_63_W0_clk),
    .W0_data(mem_0_63_W0_data),
    .W0_en(mem_0_63_W0_en),
    .W0_mask(mem_0_63_W0_mask)
  );
  assign R0_data = {R0_data_0_63,_GEN_61};
  assign mem_0_0_R0_addr = R0_addr;
  assign mem_0_0_R0_clk = R0_clk;
  assign mem_0_0_R0_en = R0_en;
  assign mem_0_0_W0_addr = W0_addr;
  assign mem_0_0_W0_clk = W0_clk;
  assign mem_0_0_W0_data = W0_data[7:0];
  assign mem_0_0_W0_en = W0_en;
  assign mem_0_0_W0_mask = W0_mask[0];
  assign mem_0_1_R0_addr = R0_addr;
  assign mem_0_1_R0_clk = R0_clk;
  assign mem_0_1_R0_en = R0_en;
  assign mem_0_1_W0_addr = W0_addr;
  assign mem_0_1_W0_clk = W0_clk;
  assign mem_0_1_W0_data = W0_data[15:8];
  assign mem_0_1_W0_en = W0_en;
  assign mem_0_1_W0_mask = W0_mask[1];
  assign mem_0_2_R0_addr = R0_addr;
  assign mem_0_2_R0_clk = R0_clk;
  assign mem_0_2_R0_en = R0_en;
  assign mem_0_2_W0_addr = W0_addr;
  assign mem_0_2_W0_clk = W0_clk;
  assign mem_0_2_W0_data = W0_data[23:16];
  assign mem_0_2_W0_en = W0_en;
  assign mem_0_2_W0_mask = W0_mask[2];
  assign mem_0_3_R0_addr = R0_addr;
  assign mem_0_3_R0_clk = R0_clk;
  assign mem_0_3_R0_en = R0_en;
  assign mem_0_3_W0_addr = W0_addr;
  assign mem_0_3_W0_clk = W0_clk;
  assign mem_0_3_W0_data = W0_data[31:24];
  assign mem_0_3_W0_en = W0_en;
  assign mem_0_3_W0_mask = W0_mask[3];
  assign mem_0_4_R0_addr = R0_addr;
  assign mem_0_4_R0_clk = R0_clk;
  assign mem_0_4_R0_en = R0_en;
  assign mem_0_4_W0_addr = W0_addr;
  assign mem_0_4_W0_clk = W0_clk;
  assign mem_0_4_W0_data = W0_data[39:32];
  assign mem_0_4_W0_en = W0_en;
  assign mem_0_4_W0_mask = W0_mask[4];
  assign mem_0_5_R0_addr = R0_addr;
  assign mem_0_5_R0_clk = R0_clk;
  assign mem_0_5_R0_en = R0_en;
  assign mem_0_5_W0_addr = W0_addr;
  assign mem_0_5_W0_clk = W0_clk;
  assign mem_0_5_W0_data = W0_data[47:40];
  assign mem_0_5_W0_en = W0_en;
  assign mem_0_5_W0_mask = W0_mask[5];
  assign mem_0_6_R0_addr = R0_addr;
  assign mem_0_6_R0_clk = R0_clk;
  assign mem_0_6_R0_en = R0_en;
  assign mem_0_6_W0_addr = W0_addr;
  assign mem_0_6_W0_clk = W0_clk;
  assign mem_0_6_W0_data = W0_data[55:48];
  assign mem_0_6_W0_en = W0_en;
  assign mem_0_6_W0_mask = W0_mask[6];
  assign mem_0_7_R0_addr = R0_addr;
  assign mem_0_7_R0_clk = R0_clk;
  assign mem_0_7_R0_en = R0_en;
  assign mem_0_7_W0_addr = W0_addr;
  assign mem_0_7_W0_clk = W0_clk;
  assign mem_0_7_W0_data = W0_data[63:56];
  assign mem_0_7_W0_en = W0_en;
  assign mem_0_7_W0_mask = W0_mask[7];
  assign mem_0_8_R0_addr = R0_addr;
  assign mem_0_8_R0_clk = R0_clk;
  assign mem_0_8_R0_en = R0_en;
  assign mem_0_8_W0_addr = W0_addr;
  assign mem_0_8_W0_clk = W0_clk;
  assign mem_0_8_W0_data = W0_data[71:64];
  assign mem_0_8_W0_en = W0_en;
  assign mem_0_8_W0_mask = W0_mask[8];
  assign mem_0_9_R0_addr = R0_addr;
  assign mem_0_9_R0_clk = R0_clk;
  assign mem_0_9_R0_en = R0_en;
  assign mem_0_9_W0_addr = W0_addr;
  assign mem_0_9_W0_clk = W0_clk;
  assign mem_0_9_W0_data = W0_data[79:72];
  assign mem_0_9_W0_en = W0_en;
  assign mem_0_9_W0_mask = W0_mask[9];
  assign mem_0_10_R0_addr = R0_addr;
  assign mem_0_10_R0_clk = R0_clk;
  assign mem_0_10_R0_en = R0_en;
  assign mem_0_10_W0_addr = W0_addr;
  assign mem_0_10_W0_clk = W0_clk;
  assign mem_0_10_W0_data = W0_data[87:80];
  assign mem_0_10_W0_en = W0_en;
  assign mem_0_10_W0_mask = W0_mask[10];
  assign mem_0_11_R0_addr = R0_addr;
  assign mem_0_11_R0_clk = R0_clk;
  assign mem_0_11_R0_en = R0_en;
  assign mem_0_11_W0_addr = W0_addr;
  assign mem_0_11_W0_clk = W0_clk;
  assign mem_0_11_W0_data = W0_data[95:88];
  assign mem_0_11_W0_en = W0_en;
  assign mem_0_11_W0_mask = W0_mask[11];
  assign mem_0_12_R0_addr = R0_addr;
  assign mem_0_12_R0_clk = R0_clk;
  assign mem_0_12_R0_en = R0_en;
  assign mem_0_12_W0_addr = W0_addr;
  assign mem_0_12_W0_clk = W0_clk;
  assign mem_0_12_W0_data = W0_data[103:96];
  assign mem_0_12_W0_en = W0_en;
  assign mem_0_12_W0_mask = W0_mask[12];
  assign mem_0_13_R0_addr = R0_addr;
  assign mem_0_13_R0_clk = R0_clk;
  assign mem_0_13_R0_en = R0_en;
  assign mem_0_13_W0_addr = W0_addr;
  assign mem_0_13_W0_clk = W0_clk;
  assign mem_0_13_W0_data = W0_data[111:104];
  assign mem_0_13_W0_en = W0_en;
  assign mem_0_13_W0_mask = W0_mask[13];
  assign mem_0_14_R0_addr = R0_addr;
  assign mem_0_14_R0_clk = R0_clk;
  assign mem_0_14_R0_en = R0_en;
  assign mem_0_14_W0_addr = W0_addr;
  assign mem_0_14_W0_clk = W0_clk;
  assign mem_0_14_W0_data = W0_data[119:112];
  assign mem_0_14_W0_en = W0_en;
  assign mem_0_14_W0_mask = W0_mask[14];
  assign mem_0_15_R0_addr = R0_addr;
  assign mem_0_15_R0_clk = R0_clk;
  assign mem_0_15_R0_en = R0_en;
  assign mem_0_15_W0_addr = W0_addr;
  assign mem_0_15_W0_clk = W0_clk;
  assign mem_0_15_W0_data = W0_data[127:120];
  assign mem_0_15_W0_en = W0_en;
  assign mem_0_15_W0_mask = W0_mask[15];
  assign mem_0_16_R0_addr = R0_addr;
  assign mem_0_16_R0_clk = R0_clk;
  assign mem_0_16_R0_en = R0_en;
  assign mem_0_16_W0_addr = W0_addr;
  assign mem_0_16_W0_clk = W0_clk;
  assign mem_0_16_W0_data = W0_data[135:128];
  assign mem_0_16_W0_en = W0_en;
  assign mem_0_16_W0_mask = W0_mask[16];
  assign mem_0_17_R0_addr = R0_addr;
  assign mem_0_17_R0_clk = R0_clk;
  assign mem_0_17_R0_en = R0_en;
  assign mem_0_17_W0_addr = W0_addr;
  assign mem_0_17_W0_clk = W0_clk;
  assign mem_0_17_W0_data = W0_data[143:136];
  assign mem_0_17_W0_en = W0_en;
  assign mem_0_17_W0_mask = W0_mask[17];
  assign mem_0_18_R0_addr = R0_addr;
  assign mem_0_18_R0_clk = R0_clk;
  assign mem_0_18_R0_en = R0_en;
  assign mem_0_18_W0_addr = W0_addr;
  assign mem_0_18_W0_clk = W0_clk;
  assign mem_0_18_W0_data = W0_data[151:144];
  assign mem_0_18_W0_en = W0_en;
  assign mem_0_18_W0_mask = W0_mask[18];
  assign mem_0_19_R0_addr = R0_addr;
  assign mem_0_19_R0_clk = R0_clk;
  assign mem_0_19_R0_en = R0_en;
  assign mem_0_19_W0_addr = W0_addr;
  assign mem_0_19_W0_clk = W0_clk;
  assign mem_0_19_W0_data = W0_data[159:152];
  assign mem_0_19_W0_en = W0_en;
  assign mem_0_19_W0_mask = W0_mask[19];
  assign mem_0_20_R0_addr = R0_addr;
  assign mem_0_20_R0_clk = R0_clk;
  assign mem_0_20_R0_en = R0_en;
  assign mem_0_20_W0_addr = W0_addr;
  assign mem_0_20_W0_clk = W0_clk;
  assign mem_0_20_W0_data = W0_data[167:160];
  assign mem_0_20_W0_en = W0_en;
  assign mem_0_20_W0_mask = W0_mask[20];
  assign mem_0_21_R0_addr = R0_addr;
  assign mem_0_21_R0_clk = R0_clk;
  assign mem_0_21_R0_en = R0_en;
  assign mem_0_21_W0_addr = W0_addr;
  assign mem_0_21_W0_clk = W0_clk;
  assign mem_0_21_W0_data = W0_data[175:168];
  assign mem_0_21_W0_en = W0_en;
  assign mem_0_21_W0_mask = W0_mask[21];
  assign mem_0_22_R0_addr = R0_addr;
  assign mem_0_22_R0_clk = R0_clk;
  assign mem_0_22_R0_en = R0_en;
  assign mem_0_22_W0_addr = W0_addr;
  assign mem_0_22_W0_clk = W0_clk;
  assign mem_0_22_W0_data = W0_data[183:176];
  assign mem_0_22_W0_en = W0_en;
  assign mem_0_22_W0_mask = W0_mask[22];
  assign mem_0_23_R0_addr = R0_addr;
  assign mem_0_23_R0_clk = R0_clk;
  assign mem_0_23_R0_en = R0_en;
  assign mem_0_23_W0_addr = W0_addr;
  assign mem_0_23_W0_clk = W0_clk;
  assign mem_0_23_W0_data = W0_data[191:184];
  assign mem_0_23_W0_en = W0_en;
  assign mem_0_23_W0_mask = W0_mask[23];
  assign mem_0_24_R0_addr = R0_addr;
  assign mem_0_24_R0_clk = R0_clk;
  assign mem_0_24_R0_en = R0_en;
  assign mem_0_24_W0_addr = W0_addr;
  assign mem_0_24_W0_clk = W0_clk;
  assign mem_0_24_W0_data = W0_data[199:192];
  assign mem_0_24_W0_en = W0_en;
  assign mem_0_24_W0_mask = W0_mask[24];
  assign mem_0_25_R0_addr = R0_addr;
  assign mem_0_25_R0_clk = R0_clk;
  assign mem_0_25_R0_en = R0_en;
  assign mem_0_25_W0_addr = W0_addr;
  assign mem_0_25_W0_clk = W0_clk;
  assign mem_0_25_W0_data = W0_data[207:200];
  assign mem_0_25_W0_en = W0_en;
  assign mem_0_25_W0_mask = W0_mask[25];
  assign mem_0_26_R0_addr = R0_addr;
  assign mem_0_26_R0_clk = R0_clk;
  assign mem_0_26_R0_en = R0_en;
  assign mem_0_26_W0_addr = W0_addr;
  assign mem_0_26_W0_clk = W0_clk;
  assign mem_0_26_W0_data = W0_data[215:208];
  assign mem_0_26_W0_en = W0_en;
  assign mem_0_26_W0_mask = W0_mask[26];
  assign mem_0_27_R0_addr = R0_addr;
  assign mem_0_27_R0_clk = R0_clk;
  assign mem_0_27_R0_en = R0_en;
  assign mem_0_27_W0_addr = W0_addr;
  assign mem_0_27_W0_clk = W0_clk;
  assign mem_0_27_W0_data = W0_data[223:216];
  assign mem_0_27_W0_en = W0_en;
  assign mem_0_27_W0_mask = W0_mask[27];
  assign mem_0_28_R0_addr = R0_addr;
  assign mem_0_28_R0_clk = R0_clk;
  assign mem_0_28_R0_en = R0_en;
  assign mem_0_28_W0_addr = W0_addr;
  assign mem_0_28_W0_clk = W0_clk;
  assign mem_0_28_W0_data = W0_data[231:224];
  assign mem_0_28_W0_en = W0_en;
  assign mem_0_28_W0_mask = W0_mask[28];
  assign mem_0_29_R0_addr = R0_addr;
  assign mem_0_29_R0_clk = R0_clk;
  assign mem_0_29_R0_en = R0_en;
  assign mem_0_29_W0_addr = W0_addr;
  assign mem_0_29_W0_clk = W0_clk;
  assign mem_0_29_W0_data = W0_data[239:232];
  assign mem_0_29_W0_en = W0_en;
  assign mem_0_29_W0_mask = W0_mask[29];
  assign mem_0_30_R0_addr = R0_addr;
  assign mem_0_30_R0_clk = R0_clk;
  assign mem_0_30_R0_en = R0_en;
  assign mem_0_30_W0_addr = W0_addr;
  assign mem_0_30_W0_clk = W0_clk;
  assign mem_0_30_W0_data = W0_data[247:240];
  assign mem_0_30_W0_en = W0_en;
  assign mem_0_30_W0_mask = W0_mask[30];
  assign mem_0_31_R0_addr = R0_addr;
  assign mem_0_31_R0_clk = R0_clk;
  assign mem_0_31_R0_en = R0_en;
  assign mem_0_31_W0_addr = W0_addr;
  assign mem_0_31_W0_clk = W0_clk;
  assign mem_0_31_W0_data = W0_data[255:248];
  assign mem_0_31_W0_en = W0_en;
  assign mem_0_31_W0_mask = W0_mask[31];
  assign mem_0_32_R0_addr = R0_addr;
  assign mem_0_32_R0_clk = R0_clk;
  assign mem_0_32_R0_en = R0_en;
  assign mem_0_32_W0_addr = W0_addr;
  assign mem_0_32_W0_clk = W0_clk;
  assign mem_0_32_W0_data = W0_data[263:256];
  assign mem_0_32_W0_en = W0_en;
  assign mem_0_32_W0_mask = W0_mask[32];
  assign mem_0_33_R0_addr = R0_addr;
  assign mem_0_33_R0_clk = R0_clk;
  assign mem_0_33_R0_en = R0_en;
  assign mem_0_33_W0_addr = W0_addr;
  assign mem_0_33_W0_clk = W0_clk;
  assign mem_0_33_W0_data = W0_data[271:264];
  assign mem_0_33_W0_en = W0_en;
  assign mem_0_33_W0_mask = W0_mask[33];
  assign mem_0_34_R0_addr = R0_addr;
  assign mem_0_34_R0_clk = R0_clk;
  assign mem_0_34_R0_en = R0_en;
  assign mem_0_34_W0_addr = W0_addr;
  assign mem_0_34_W0_clk = W0_clk;
  assign mem_0_34_W0_data = W0_data[279:272];
  assign mem_0_34_W0_en = W0_en;
  assign mem_0_34_W0_mask = W0_mask[34];
  assign mem_0_35_R0_addr = R0_addr;
  assign mem_0_35_R0_clk = R0_clk;
  assign mem_0_35_R0_en = R0_en;
  assign mem_0_35_W0_addr = W0_addr;
  assign mem_0_35_W0_clk = W0_clk;
  assign mem_0_35_W0_data = W0_data[287:280];
  assign mem_0_35_W0_en = W0_en;
  assign mem_0_35_W0_mask = W0_mask[35];
  assign mem_0_36_R0_addr = R0_addr;
  assign mem_0_36_R0_clk = R0_clk;
  assign mem_0_36_R0_en = R0_en;
  assign mem_0_36_W0_addr = W0_addr;
  assign mem_0_36_W0_clk = W0_clk;
  assign mem_0_36_W0_data = W0_data[295:288];
  assign mem_0_36_W0_en = W0_en;
  assign mem_0_36_W0_mask = W0_mask[36];
  assign mem_0_37_R0_addr = R0_addr;
  assign mem_0_37_R0_clk = R0_clk;
  assign mem_0_37_R0_en = R0_en;
  assign mem_0_37_W0_addr = W0_addr;
  assign mem_0_37_W0_clk = W0_clk;
  assign mem_0_37_W0_data = W0_data[303:296];
  assign mem_0_37_W0_en = W0_en;
  assign mem_0_37_W0_mask = W0_mask[37];
  assign mem_0_38_R0_addr = R0_addr;
  assign mem_0_38_R0_clk = R0_clk;
  assign mem_0_38_R0_en = R0_en;
  assign mem_0_38_W0_addr = W0_addr;
  assign mem_0_38_W0_clk = W0_clk;
  assign mem_0_38_W0_data = W0_data[311:304];
  assign mem_0_38_W0_en = W0_en;
  assign mem_0_38_W0_mask = W0_mask[38];
  assign mem_0_39_R0_addr = R0_addr;
  assign mem_0_39_R0_clk = R0_clk;
  assign mem_0_39_R0_en = R0_en;
  assign mem_0_39_W0_addr = W0_addr;
  assign mem_0_39_W0_clk = W0_clk;
  assign mem_0_39_W0_data = W0_data[319:312];
  assign mem_0_39_W0_en = W0_en;
  assign mem_0_39_W0_mask = W0_mask[39];
  assign mem_0_40_R0_addr = R0_addr;
  assign mem_0_40_R0_clk = R0_clk;
  assign mem_0_40_R0_en = R0_en;
  assign mem_0_40_W0_addr = W0_addr;
  assign mem_0_40_W0_clk = W0_clk;
  assign mem_0_40_W0_data = W0_data[327:320];
  assign mem_0_40_W0_en = W0_en;
  assign mem_0_40_W0_mask = W0_mask[40];
  assign mem_0_41_R0_addr = R0_addr;
  assign mem_0_41_R0_clk = R0_clk;
  assign mem_0_41_R0_en = R0_en;
  assign mem_0_41_W0_addr = W0_addr;
  assign mem_0_41_W0_clk = W0_clk;
  assign mem_0_41_W0_data = W0_data[335:328];
  assign mem_0_41_W0_en = W0_en;
  assign mem_0_41_W0_mask = W0_mask[41];
  assign mem_0_42_R0_addr = R0_addr;
  assign mem_0_42_R0_clk = R0_clk;
  assign mem_0_42_R0_en = R0_en;
  assign mem_0_42_W0_addr = W0_addr;
  assign mem_0_42_W0_clk = W0_clk;
  assign mem_0_42_W0_data = W0_data[343:336];
  assign mem_0_42_W0_en = W0_en;
  assign mem_0_42_W0_mask = W0_mask[42];
  assign mem_0_43_R0_addr = R0_addr;
  assign mem_0_43_R0_clk = R0_clk;
  assign mem_0_43_R0_en = R0_en;
  assign mem_0_43_W0_addr = W0_addr;
  assign mem_0_43_W0_clk = W0_clk;
  assign mem_0_43_W0_data = W0_data[351:344];
  assign mem_0_43_W0_en = W0_en;
  assign mem_0_43_W0_mask = W0_mask[43];
  assign mem_0_44_R0_addr = R0_addr;
  assign mem_0_44_R0_clk = R0_clk;
  assign mem_0_44_R0_en = R0_en;
  assign mem_0_44_W0_addr = W0_addr;
  assign mem_0_44_W0_clk = W0_clk;
  assign mem_0_44_W0_data = W0_data[359:352];
  assign mem_0_44_W0_en = W0_en;
  assign mem_0_44_W0_mask = W0_mask[44];
  assign mem_0_45_R0_addr = R0_addr;
  assign mem_0_45_R0_clk = R0_clk;
  assign mem_0_45_R0_en = R0_en;
  assign mem_0_45_W0_addr = W0_addr;
  assign mem_0_45_W0_clk = W0_clk;
  assign mem_0_45_W0_data = W0_data[367:360];
  assign mem_0_45_W0_en = W0_en;
  assign mem_0_45_W0_mask = W0_mask[45];
  assign mem_0_46_R0_addr = R0_addr;
  assign mem_0_46_R0_clk = R0_clk;
  assign mem_0_46_R0_en = R0_en;
  assign mem_0_46_W0_addr = W0_addr;
  assign mem_0_46_W0_clk = W0_clk;
  assign mem_0_46_W0_data = W0_data[375:368];
  assign mem_0_46_W0_en = W0_en;
  assign mem_0_46_W0_mask = W0_mask[46];
  assign mem_0_47_R0_addr = R0_addr;
  assign mem_0_47_R0_clk = R0_clk;
  assign mem_0_47_R0_en = R0_en;
  assign mem_0_47_W0_addr = W0_addr;
  assign mem_0_47_W0_clk = W0_clk;
  assign mem_0_47_W0_data = W0_data[383:376];
  assign mem_0_47_W0_en = W0_en;
  assign mem_0_47_W0_mask = W0_mask[47];
  assign mem_0_48_R0_addr = R0_addr;
  assign mem_0_48_R0_clk = R0_clk;
  assign mem_0_48_R0_en = R0_en;
  assign mem_0_48_W0_addr = W0_addr;
  assign mem_0_48_W0_clk = W0_clk;
  assign mem_0_48_W0_data = W0_data[391:384];
  assign mem_0_48_W0_en = W0_en;
  assign mem_0_48_W0_mask = W0_mask[48];
  assign mem_0_49_R0_addr = R0_addr;
  assign mem_0_49_R0_clk = R0_clk;
  assign mem_0_49_R0_en = R0_en;
  assign mem_0_49_W0_addr = W0_addr;
  assign mem_0_49_W0_clk = W0_clk;
  assign mem_0_49_W0_data = W0_data[399:392];
  assign mem_0_49_W0_en = W0_en;
  assign mem_0_49_W0_mask = W0_mask[49];
  assign mem_0_50_R0_addr = R0_addr;
  assign mem_0_50_R0_clk = R0_clk;
  assign mem_0_50_R0_en = R0_en;
  assign mem_0_50_W0_addr = W0_addr;
  assign mem_0_50_W0_clk = W0_clk;
  assign mem_0_50_W0_data = W0_data[407:400];
  assign mem_0_50_W0_en = W0_en;
  assign mem_0_50_W0_mask = W0_mask[50];
  assign mem_0_51_R0_addr = R0_addr;
  assign mem_0_51_R0_clk = R0_clk;
  assign mem_0_51_R0_en = R0_en;
  assign mem_0_51_W0_addr = W0_addr;
  assign mem_0_51_W0_clk = W0_clk;
  assign mem_0_51_W0_data = W0_data[415:408];
  assign mem_0_51_W0_en = W0_en;
  assign mem_0_51_W0_mask = W0_mask[51];
  assign mem_0_52_R0_addr = R0_addr;
  assign mem_0_52_R0_clk = R0_clk;
  assign mem_0_52_R0_en = R0_en;
  assign mem_0_52_W0_addr = W0_addr;
  assign mem_0_52_W0_clk = W0_clk;
  assign mem_0_52_W0_data = W0_data[423:416];
  assign mem_0_52_W0_en = W0_en;
  assign mem_0_52_W0_mask = W0_mask[52];
  assign mem_0_53_R0_addr = R0_addr;
  assign mem_0_53_R0_clk = R0_clk;
  assign mem_0_53_R0_en = R0_en;
  assign mem_0_53_W0_addr = W0_addr;
  assign mem_0_53_W0_clk = W0_clk;
  assign mem_0_53_W0_data = W0_data[431:424];
  assign mem_0_53_W0_en = W0_en;
  assign mem_0_53_W0_mask = W0_mask[53];
  assign mem_0_54_R0_addr = R0_addr;
  assign mem_0_54_R0_clk = R0_clk;
  assign mem_0_54_R0_en = R0_en;
  assign mem_0_54_W0_addr = W0_addr;
  assign mem_0_54_W0_clk = W0_clk;
  assign mem_0_54_W0_data = W0_data[439:432];
  assign mem_0_54_W0_en = W0_en;
  assign mem_0_54_W0_mask = W0_mask[54];
  assign mem_0_55_R0_addr = R0_addr;
  assign mem_0_55_R0_clk = R0_clk;
  assign mem_0_55_R0_en = R0_en;
  assign mem_0_55_W0_addr = W0_addr;
  assign mem_0_55_W0_clk = W0_clk;
  assign mem_0_55_W0_data = W0_data[447:440];
  assign mem_0_55_W0_en = W0_en;
  assign mem_0_55_W0_mask = W0_mask[55];
  assign mem_0_56_R0_addr = R0_addr;
  assign mem_0_56_R0_clk = R0_clk;
  assign mem_0_56_R0_en = R0_en;
  assign mem_0_56_W0_addr = W0_addr;
  assign mem_0_56_W0_clk = W0_clk;
  assign mem_0_56_W0_data = W0_data[455:448];
  assign mem_0_56_W0_en = W0_en;
  assign mem_0_56_W0_mask = W0_mask[56];
  assign mem_0_57_R0_addr = R0_addr;
  assign mem_0_57_R0_clk = R0_clk;
  assign mem_0_57_R0_en = R0_en;
  assign mem_0_57_W0_addr = W0_addr;
  assign mem_0_57_W0_clk = W0_clk;
  assign mem_0_57_W0_data = W0_data[463:456];
  assign mem_0_57_W0_en = W0_en;
  assign mem_0_57_W0_mask = W0_mask[57];
  assign mem_0_58_R0_addr = R0_addr;
  assign mem_0_58_R0_clk = R0_clk;
  assign mem_0_58_R0_en = R0_en;
  assign mem_0_58_W0_addr = W0_addr;
  assign mem_0_58_W0_clk = W0_clk;
  assign mem_0_58_W0_data = W0_data[471:464];
  assign mem_0_58_W0_en = W0_en;
  assign mem_0_58_W0_mask = W0_mask[58];
  assign mem_0_59_R0_addr = R0_addr;
  assign mem_0_59_R0_clk = R0_clk;
  assign mem_0_59_R0_en = R0_en;
  assign mem_0_59_W0_addr = W0_addr;
  assign mem_0_59_W0_clk = W0_clk;
  assign mem_0_59_W0_data = W0_data[479:472];
  assign mem_0_59_W0_en = W0_en;
  assign mem_0_59_W0_mask = W0_mask[59];
  assign mem_0_60_R0_addr = R0_addr;
  assign mem_0_60_R0_clk = R0_clk;
  assign mem_0_60_R0_en = R0_en;
  assign mem_0_60_W0_addr = W0_addr;
  assign mem_0_60_W0_clk = W0_clk;
  assign mem_0_60_W0_data = W0_data[487:480];
  assign mem_0_60_W0_en = W0_en;
  assign mem_0_60_W0_mask = W0_mask[60];
  assign mem_0_61_R0_addr = R0_addr;
  assign mem_0_61_R0_clk = R0_clk;
  assign mem_0_61_R0_en = R0_en;
  assign mem_0_61_W0_addr = W0_addr;
  assign mem_0_61_W0_clk = W0_clk;
  assign mem_0_61_W0_data = W0_data[495:488];
  assign mem_0_61_W0_en = W0_en;
  assign mem_0_61_W0_mask = W0_mask[61];
  assign mem_0_62_R0_addr = R0_addr;
  assign mem_0_62_R0_clk = R0_clk;
  assign mem_0_62_R0_en = R0_en;
  assign mem_0_62_W0_addr = W0_addr;
  assign mem_0_62_W0_clk = W0_clk;
  assign mem_0_62_W0_data = W0_data[503:496];
  assign mem_0_62_W0_en = W0_en;
  assign mem_0_62_W0_mask = W0_mask[62];
  assign mem_0_63_R0_addr = R0_addr;
  assign mem_0_63_R0_clk = R0_clk;
  assign mem_0_63_R0_en = R0_en;
  assign mem_0_63_W0_addr = W0_addr;
  assign mem_0_63_W0_clk = W0_clk;
  assign mem_0_63_W0_data = W0_data[511:504];
  assign mem_0_63_W0_en = W0_en;
  assign mem_0_63_W0_mask = W0_mask[63];
endmodule
module tag_array_0_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [83:0] RW0_wdata,
  output [83:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input  [3:0]  RW0_wmask
);
  wire [5:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [20:0] mem_0_0_RW0_wdata;
  wire [20:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [5:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [20:0] mem_0_1_RW0_wdata;
  wire [20:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [5:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [20:0] mem_0_2_RW0_wdata;
  wire [20:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [5:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [20:0] mem_0_3_RW0_wdata;
  wire [20:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [20:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [20:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [20:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [20:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [41:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [62:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [83:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [41:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [62:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  split_tag_array_0_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[20:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[41:21];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[62:42];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[83:63];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
endmodule
module data_arrays_0_0_ext(
  input  [7:0]   RW0_addr,
  input          RW0_clk,
  input  [127:0] RW0_wdata,
  output [127:0] RW0_rdata,
  input          RW0_en,
  input          RW0_wmode,
  input  [3:0]   RW0_wmask
);
  wire [7:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [31:0] mem_0_0_RW0_wdata;
  wire [31:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [7:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [31:0] mem_0_1_RW0_wdata;
  wire [31:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [7:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [31:0] mem_0_2_RW0_wdata;
  wire [31:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [7:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [31:0] mem_0_3_RW0_wdata;
  wire [31:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [31:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [31:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [31:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [31:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [63:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [95:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [127:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [63:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [95:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  split_data_arrays_0_0_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[31:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[63:32];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[95:64];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[127:96];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask[3];
endmodule
module l2_tlb_ram_0_ext(
  input  [8:0]  RW0_addr,
  input         RW0_clk,
  input  [44:0] RW0_wdata,
  output [44:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
  wire [8:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [44:0] mem_0_0_RW0_wdata;
  wire [44:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire [44:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [44:0] RW0_rdata_0 = RW0_rdata_0_0;
  split_l2_tlb_ram_0_ext mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata = mem_0_0_RW0_rdata;
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata;
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
endmodule
module split_cc_dir_ext(
  input  [9:0]  RW0_addr,
  input         RW0_clk,
  input  [15:0] RW0_wdata,
  output [15:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ram [0:1023];
  wire  ram_RW_0_r_en;
  wire [9:0] ram_RW_0_r_addr;
  wire [15:0] ram_RW_0_r_data;
  wire [15:0] ram_RW_0_w_data;
  wire [9:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [9:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_cc_banks_0_ext(
  input  [12:0] RW0_addr,
  input         RW0_clk,
  input  [63:0] RW0_wdata,
  output [63:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:8191];
  wire  ram_RW_0_r_en;
  wire [12:0] ram_RW_0_r_addr;
  wire [63:0] ram_RW_0_r_data;
  wire [63:0] ram_RW_0_w_data;
  wire [12:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [12:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[12:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_data_arrays_0_ext(
  input  [7:0] RW0_addr,
  input        RW0_clk,
  input  [7:0] RW0_wdata,
  output [7:0] RW0_rdata,
  input        RW0_en,
  input        RW0_wmode,
  input        RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:255];
  wire  ram_RW_0_r_en;
  wire [7:0] ram_RW_0_r_addr;
  wire [7:0] ram_RW_0_r_data;
  wire [7:0] ram_RW_0_w_data;
  wire [7:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [7:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_tag_array_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [21:0] RW0_wdata,
  output [21:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [21:0] ram [0:63];
  wire  ram_RW_0_r_en;
  wire [5:0] ram_RW_0_r_addr;
  wire [21:0] ram_RW_0_r_data;
  wire [21:0] ram_RW_0_w_data;
  wire [5:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[21:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_mem_ext(
  input  [11:0] RW0_addr,
  input         RW0_clk,
  input  [7:0]  RW0_wdata,
  output [7:0]  RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:4095];
  wire  ram_RW_0_r_en;
  wire [11:0] ram_RW_0_r_addr;
  wire [7:0] ram_RW_0_r_data;
  wire [7:0] ram_RW_0_w_data;
  wire [11:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [11:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_mem_0_ext(
  input  [8:0] R0_addr,
  input        R0_clk,
  output [7:0] R0_data,
  input        R0_en,
  input  [8:0] W0_addr,
  input        W0_clk,
  input  [7:0] W0_data,
  input        W0_en,
  input        W0_mask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:511];
  wire  ram_R_0_en;
  wire [8:0] ram_R_0_addr;
  wire [7:0] ram_R_0_data;
  wire [7:0] ram_W_0_data;
  wire [8:0] ram_W_0_addr;
  wire  ram_W_0_mask;
  wire  ram_W_0_en;
  reg  ram_R_0_en_pipe_0;
  reg [8:0] ram_R_0_addr_pipe_0;
  assign ram_R_0_en = ram_R_0_en_pipe_0;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr];
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data;
  always @(posedge W0_clk) begin
    if (ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data;
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_tag_array_0_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [20:0] RW0_wdata,
  output [20:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] ram [0:63];
  wire  ram_RW_0_r_en;
  wire [5:0] ram_RW_0_r_addr;
  wire [20:0] ram_RW_0_r_data;
  wire [20:0] ram_RW_0_w_data;
  wire [5:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[20:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_data_arrays_0_0_ext(
  input  [7:0]  RW0_addr,
  input         RW0_clk,
  input  [31:0] RW0_wdata,
  output [31:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram [0:255];
  wire  ram_RW_0_r_en;
  wire [7:0] ram_RW_0_r_addr;
  wire [31:0] ram_RW_0_r_data;
  wire [31:0] ram_RW_0_w_data;
  wire [7:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [7:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module split_l2_tlb_ram_0_ext(
  input  [8:0]  RW0_addr,
  input         RW0_clk,
  input  [44:0] RW0_wdata,
  output [44:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [44:0] ram [0:511];
  wire  ram_RW_0_r_en;
  wire [8:0] ram_RW_0_r_addr;
  wire [44:0] ram_RW_0_r_data;
  wire [44:0] ram_RW_0_w_data;
  wire [8:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [8:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    ram[initvar] = _RAND_0[44:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
